* NGSPICE file created from heichips25_CORDIC.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

.subckt heichips25_CORDIC VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
X_6914_ net270 VGND VPWR _0509_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[8\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_1
X_6845_ net580 VGND VPWR _0454_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[2\]
+ clknet_leaf_65_clk sg13g2_dfrbpq_2
X_6776_ net649 VGND VPWR net1328 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[9\]
+ clknet_leaf_58_clk sg13g2_dfrbpq_1
XFILLER_22_166 VPWR VGND sg13g2_fill_1
X_6871__343 VPWR VGND net343 sg13g2_tiehi
X_3988_ _0989_ net449 _0987_ VPWR VGND sg13g2_nand2b_1
X_5727_ VGND VPWR _2415_ _2419_ _2422_ _2417_ sg13g2_a21oi_1
X_5658_ _2356_ _2361_ _2362_ VPWR VGND sg13g2_nor2_1
X_4609_ _1494_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[9\] _1493_
+ VPWR VGND sg13g2_xnor2_1
X_5589_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[5\] _2302_ _2303_
+ VPWR VGND sg13g2_and2_1
Xhold362 _0362_ VPWR VGND net1119 sg13g2_dlygate4sd3_1
Xhold351 _2909_ VPWR VGND net1108 sg13g2_dlygate4sd3_1
Xhold340 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[1\] VPWR VGND net1097
+ sg13g2_dlygate4sd3_1
Xhold373 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[11\] VPWR VGND net1130
+ sg13g2_dlygate4sd3_1
Xhold395 _0091_ VPWR VGND net1152 sg13g2_dlygate4sd3_1
Xhold384 _0128_ VPWR VGND net1141 sg13g2_dlygate4sd3_1
XFILLER_26_52 VPWR VGND sg13g2_fill_1
XFILLER_27_995 VPWR VGND sg13g2_decap_8
XFILLER_6_811 VPWR VGND sg13g2_decap_8
XFILLER_10_873 VPWR VGND sg13g2_decap_8
XFILLER_6_888 VPWR VGND sg13g2_decap_8
XFILLER_47_8 VPWR VGND sg13g2_decap_8
XFILLER_3_1018 VPWR VGND sg13g2_decap_8
X_6902__553 VPWR VGND net737 sg13g2_tiehi
XFILLER_18_940 VPWR VGND sg13g2_decap_8
XFILLER_45_781 VPWR VGND sg13g2_fill_1
X_4960_ _1789_ net399 net1494 _1778_ net1464 VPWR VGND sg13g2_a22oi_1
XFILLER_33_921 VPWR VGND sg13g2_fill_1
X_4891_ net389 VPWR _1731_ VGND net1167 net1533 sg13g2_o21ai_1
X_3911_ VGND VPWR net863 _0925_ _0041_ _0926_ sg13g2_a21oi_1
X_6630_ net92 VGND VPWR _0239_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[3\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_1
X_3842_ net950 _0876_ _0877_ VPWR VGND sg13g2_nor2_1
X_6561_ net161 VGND VPWR net833 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].z_sign
+ clknet_leaf_40_clk sg13g2_dfrbpq_2
X_3773_ _0542_ net936 net950 net874 _0821_ VPWR VGND sg13g2_nor4_1
X_5512_ _2239_ net418 net1358 VPWR VGND sg13g2_nand2_1
X_6419__342 VPWR VGND net342 sg13g2_tiehi
X_6492_ net230 VGND VPWR _0101_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[6\]
+ clknet_leaf_45_clk sg13g2_dfrbpq_1
X_5443_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[1\] _2180_
+ _2182_ VPWR VGND sg13g2_nor2_1
X_5374_ VGND VPWR _2117_ _2122_ _0307_ _2123_ sg13g2_a21oi_1
X_4325_ net542 net817 _1260_ VPWR VGND sg13g2_nor2b_1
X_4256_ _1195_ VPWR _1202_ VGND net531 _0584_ sg13g2_o21ai_1
X_4187_ net437 _1143_ _1144_ _0099_ VPWR VGND sg13g2_nor3_1
XFILLER_27_236 VPWR VGND sg13g2_fill_2
X_6828_ net597 VGND VPWR _0437_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[8\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_2
X_6759_ net666 VGND VPWR net1205 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[4\]
+ clknet_leaf_30_clk sg13g2_dfrbpq_1
XFILLER_3_836 VPWR VGND sg13g2_decap_8
Xhold170 _2904_ VPWR VGND net927 sg13g2_dlygate4sd3_1
Xhold192 _0060_ VPWR VGND net949 sg13g2_dlygate4sd3_1
Xhold181 _0023_ VPWR VGND net938 sg13g2_dlygate4sd3_1
XFILLER_46_534 VPWR VGND sg13g2_fill_1
XFILLER_15_976 VPWR VGND sg13g2_decap_8
XFILLER_10_692 VPWR VGND sg13g2_fill_2
X_4110_ _1081_ net499 _1080_ VPWR VGND sg13g2_nand2_1
X_5090_ net1034 _1883_ _0262_ VPWR VGND sg13g2_nor2b_1
X_4041_ _1028_ _1032_ _0939_ _1034_ VPWR VGND _1033_ sg13g2_nand4_1
X_5992_ _2639_ net414 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[8\]
+ VPWR VGND sg13g2_nand2_1
X_4943_ net469 VPWR _1775_ VGND _1769_ _1774_ sg13g2_o21ai_1
X_6613_ net109 VGND VPWR net1342 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[11\]
+ clknet_leaf_25_clk sg13g2_dfrbpq_2
X_4874_ _1717_ net1493 _1716_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_423 VPWR VGND sg13g2_fill_2
X_3825_ _0812_ _0816_ _0864_ _0865_ VPWR VGND sg13g2_nor3_1
XFILLER_21_968 VPWR VGND sg13g2_decap_8
X_6544_ net178 VGND VPWR net1333 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[7\]
+ clknet_leaf_37_clk sg13g2_dfrbpq_1
X_3756_ _0796_ _0785_ _0795_ _0809_ VPWR VGND sg13g2_a21o_1
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk VPWR VGND sg13g2_buf_8
X_6475_ net247 VGND VPWR _0084_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[1\]
+ clknet_leaf_38_clk sg13g2_dfrbpq_1
X_5426_ _2167_ net1367 _2166_ VPWR VGND sg13g2_nand2_1
X_3687_ VPWR VGND _0733_ _0739_ _0736_ _0730_ _0740_ _0734_ sg13g2_a221oi_1
X_5357_ VGND VPWR _2103_ _2107_ _0305_ _2108_ sg13g2_a21oi_1
X_4308_ _1241_ _1242_ _1247_ VPWR VGND sg13g2_nor2_1
X_5288_ VGND VPWR _2051_ _2050_ _2048_ sg13g2_or2_1
X_4239_ net479 VPWR _1188_ VGND net962 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[0\]
+ sg13g2_o21ai_1
XFILLER_28_589 VPWR VGND sg13g2_fill_2
XFILLER_43_559 VPWR VGND sg13g2_fill_2
XFILLER_12_935 VPWR VGND sg13g2_decap_8
XFILLER_23_261 VPWR VGND sg13g2_fill_2
XFILLER_7_405 VPWR VGND sg13g2_fill_1
XFILLER_3_611 VPWR VGND sg13g2_fill_1
Xfanout480 net491 net480 VPWR VGND sg13g2_buf_8
Xfanout491 net505 net491 VPWR VGND sg13g2_buf_8
X_4590_ _1480_ _0608_ net1086 VPWR VGND sg13g2_nand2_1
X_3610_ VGND VPWR _0663_ _0662_ _0661_ sg13g2_or2_1
X_3541_ VPWR _0611_ net1272 VGND sg13g2_inv_1
X_3472_ VPWR _0542_ u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[6\] VGND sg13g2_inv_1
X_6260_ VGND VPWR _2860_ _2862_ _0454_ net421 sg13g2_a21oi_1
XFILLER_9_1002 VPWR VGND sg13g2_decap_8
X_5211_ _1983_ _1987_ _1989_ VPWR VGND sg13g2_and2_1
X_6191_ _2810_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[12\] _2809_
+ VPWR VGND sg13g2_xnor2_1
X_5142_ VGND VPWR net1163 _1928_ _0268_ _1930_ sg13g2_a21oi_1
X_5073_ VGND VPWR _1880_ _1881_ _0247_ _1882_ sg13g2_a21oi_1
X_4024_ _1020_ _1016_ _1019_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_397 VPWR VGND sg13g2_fill_2
X_5975_ VGND VPWR _2628_ _2629_ _0401_ _2630_ sg13g2_a21oi_1
X_4926_ VPWR _1761_ _1760_ VGND sg13g2_inv_1
X_4857_ net483 VPWR _1703_ VGND net998 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[0\]
+ sg13g2_o21ai_1
X_3808_ _0787_ _0769_ _0851_ VPWR VGND sg13g2_xor2_1
XFILLER_21_798 VPWR VGND sg13g2_fill_1
X_4788_ VGND VPWR _1645_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[10\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[9\] sg13g2_or2_1
X_6527_ net195 VGND VPWR net1453 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[3\]
+ clknet_leaf_41_clk sg13g2_dfrbpq_2
X_3739_ _0792_ _0789_ _0791_ VPWR VGND sg13g2_nand2b_1
X_6458_ net277 VGND VPWR _0067_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[11\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
X_5409_ _2152_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[5\] _2151_
+ VPWR VGND sg13g2_xnor2_1
X_6389_ VGND VPWR _2892_ _2893_ _0475_ _2890_ sg13g2_a21oi_1
XFILLER_0_647 VPWR VGND sg13g2_decap_8
XFILLER_18_53 VPWR VGND sg13g2_fill_1
XFILLER_15_1018 VPWR VGND sg13g2_decap_8
XFILLER_8_758 VPWR VGND sg13g2_fill_1
XFILLER_4_986 VPWR VGND sg13g2_decap_8
XFILLER_34_323 VPWR VGND sg13g2_fill_1
XFILLER_22_529 VPWR VGND sg13g2_fill_1
X_5760_ net517 net1084 _2448_ VPWR VGND sg13g2_nor2b_1
X_5691_ _2385_ _2390_ _2391_ VPWR VGND sg13g2_nor2_1
X_4711_ VPWR _1581_ _1580_ VGND sg13g2_inv_1
X_4642_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[12\] net537 _1515_
+ _1523_ VPWR VGND sg13g2_a21o_1
Xhold703 _0192_ VPWR VGND net1460 sg13g2_dlygate4sd3_1
X_4573_ _1466_ _1459_ _1462_ _1464_ VPWR VGND sg13g2_and3_1
Xhold736 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[10\] VPWR
+ VGND net1493 sg13g2_dlygate4sd3_1
X_3524_ VPWR _0594_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[2\]
+ VGND sg13g2_inv_1
Xhold725 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[9\] VPWR VGND net1482
+ sg13g2_dlygate4sd3_1
X_6312_ net758 net422 _0486_ VPWR VGND sg13g2_nor2_1
Xhold714 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[6\] VPWR VGND net1471
+ sg13g2_dlygate4sd3_1
Xhold747 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[9\] VPWR VGND net1504
+ sg13g2_dlygate4sd3_1
Xhold769 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[8\] VPWR VGND net1526
+ sg13g2_dlygate4sd3_1
X_6243_ _2851_ net455 _2850_ VPWR VGND sg13g2_nand2_1
Xhold758 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[7\] VPWR VGND net1515
+ sg13g2_dlygate4sd3_1
X_6174_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[10\] _2794_ _2795_
+ VPWR VGND sg13g2_nor2_1
X_5125_ _0266_ net492 _1914_ _1915_ VPWR VGND sg13g2_and3_1
X_5056_ _1869_ _1865_ _1867_ _1868_ VPWR VGND sg13g2_and3_1
X_4007_ VGND VPWR u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[2\]
+ net549 _1005_ _1001_ sg13g2_a21oi_1
XFILLER_26_824 VPWR VGND sg13g2_fill_1
XFILLER_26_835 VPWR VGND sg13g2_fill_1
X_5958_ _2616_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[12\] _2615_
+ VPWR VGND sg13g2_xnor2_1
X_6497__225 VPWR VGND net225 sg13g2_tiehi
XFILLER_41_849 VPWR VGND sg13g2_fill_2
X_4909_ VGND VPWR _1747_ _1746_ _1744_ sg13g2_or2_1
X_5889_ net512 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[2\] _2556_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_1_945 VPWR VGND sg13g2_decap_8
X_6881__323 VPWR VGND net323 sg13g2_tiehi
Xhold41 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[0\] VPWR VGND net798
+ sg13g2_dlygate4sd3_1
XFILLER_0_488 VPWR VGND sg13g2_fill_1
Xhold30 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[6\] VPWR VGND net787
+ sg13g2_dlygate4sd3_1
Xhold63 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[3\] VPWR VGND net820
+ sg13g2_dlygate4sd3_1
Xhold74 u_angle_cordic_12b_pmod.u_vga_top.clk_div_cnt\[1\] VPWR VGND net831 sg13g2_dlygate4sd3_1
Xhold52 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[0\] VPWR VGND net809
+ sg13g2_dlygate4sd3_1
Xhold85 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[8\] VPWR VGND net842 sg13g2_dlygate4sd3_1
Xhold96 _0327_ VPWR VGND net853 sg13g2_dlygate4sd3_1
XFILLER_17_835 VPWR VGND sg13g2_fill_2
XFILLER_43_120 VPWR VGND sg13g2_fill_1
XFILLER_4_783 VPWR VGND sg13g2_decap_8
X_6861_ net363 VGND VPWR _0470_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[5\]
+ clknet_leaf_63_clk sg13g2_dfrbpq_2
X_5812_ _2489_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[3\]
+ _2490_ VPWR VGND sg13g2_xor2_1
X_6858__369 VPWR VGND net369 sg13g2_tiehi
X_6792_ net633 VGND VPWR net1324 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[10\]
+ clknet_leaf_9_clk sg13g2_dfrbpq_2
X_5743_ _2434_ net412 net1280 VPWR VGND sg13g2_nand2_1
X_5674_ _2374_ net1443 _2376_ VPWR VGND sg13g2_xor2_1
X_4625_ net538 _1507_ _1508_ VPWR VGND sg13g2_nor2_1
X_4556_ _1449_ _1451_ _1447_ _1452_ VPWR VGND sg13g2_nand3_1
Xhold500 _0303_ VPWR VGND net1257 sg13g2_dlygate4sd3_1
Xhold511 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[9\] VPWR VGND net1268
+ sg13g2_dlygate4sd3_1
X_3507_ VPWR _0577_ net1554 VGND sg13g2_inv_1
Xhold533 _0271_ VPWR VGND net1290 sg13g2_dlygate4sd3_1
Xhold522 _1199_ VPWR VGND net1279 sg13g2_dlygate4sd3_1
Xhold544 _0106_ VPWR VGND net1301 sg13g2_dlygate4sd3_1
Xhold555 _0187_ VPWR VGND net1312 sg13g2_dlygate4sd3_1
Xhold577 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[8\] VPWR VGND net1334
+ sg13g2_dlygate4sd3_1
Xhold588 _0438_ VPWR VGND net1345 sg13g2_dlygate4sd3_1
Xhold566 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[10\] VPWR
+ VGND net1323 sg13g2_dlygate4sd3_1
X_4487_ _1395_ _0601_ _1394_ VPWR VGND sg13g2_xnor2_1
Xhold599 _1127_ VPWR VGND net1356 sg13g2_dlygate4sd3_1
X_6226_ _2837_ net417 net1235 VPWR VGND sg13g2_nand2_1
X_6157_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[8\] _2779_ _2780_
+ VPWR VGND sg13g2_nor2_1
X_5108_ net526 _1892_ _1900_ VPWR VGND sg13g2_nor2_1
X_6429__322 VPWR VGND net322 sg13g2_tiehi
X_6088_ _2719_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[10\] _2721_
+ VPWR VGND sg13g2_xor2_1
X_5039_ VGND VPWR _1851_ _1852_ _0241_ _1854_ sg13g2_a21oi_1
Xoutput20 net20 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_742 VPWR VGND sg13g2_decap_8
XFILLER_29_470 VPWR VGND sg13g2_fill_1
XFILLER_29_481 VPWR VGND sg13g2_fill_2
XFILLER_36_429 VPWR VGND sg13g2_fill_1
X_6640__82 VPWR VGND net82 sg13g2_tiehi
XFILLER_9_897 VPWR VGND sg13g2_decap_8
X_4410_ net1374 _1329_ _1330_ VPWR VGND sg13g2_and2_1
X_5390_ _2132_ net1479 _2137_ VPWR VGND sg13g2_xor2_1
X_4341_ _1273_ net410 net1080 VPWR VGND sg13g2_nand2_1
XFILLER_28_1006 VPWR VGND sg13g2_decap_8
X_4272_ _1215_ _1216_ _0112_ VPWR VGND sg13g2_nor2b_1
X_6011_ net1047 _2652_ _0414_ VPWR VGND sg13g2_nor2b_1
X_6487__235 VPWR VGND net235 sg13g2_tiehi
XFILLER_11_0 VPWR VGND sg13g2_fill_2
X_6913_ net272 VGND VPWR net1109 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[7\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_35_451 VPWR VGND sg13g2_fill_1
X_6844_ net581 VGND VPWR _0453_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[1\]
+ clknet_leaf_64_clk sg13g2_dfrbpq_2
X_6775_ net650 VGND VPWR _0384_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[8\]
+ clknet_leaf_58_clk sg13g2_dfrbpq_2
X_3987_ net423 _0987_ _0988_ VPWR VGND sg13g2_nor2_1
X_5726_ _2420_ _2421_ _0361_ VPWR VGND sg13g2_nor2b_1
X_6494__228 VPWR VGND net228 sg13g2_tiehi
X_5657_ _2361_ net1446 _2359_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_1010 VPWR VGND sg13g2_decap_8
X_4608_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].z_sign u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[8\]
+ _1493_ VPWR VGND sg13g2_nor2b_1
X_5588_ _2301_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[5\]
+ _2302_ VPWR VGND sg13g2_xor2_1
Xhold341 _0134_ VPWR VGND net1098 sg13g2_dlygate4sd3_1
X_4539_ VPWR _1439_ _1438_ VGND sg13g2_inv_1
Xhold352 _0508_ VPWR VGND net1109 sg13g2_dlygate4sd3_1
Xhold330 _1481_ VPWR VGND net1087 sg13g2_dlygate4sd3_1
Xhold385 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[10\] VPWR VGND net1142
+ sg13g2_dlygate4sd3_1
Xhold374 _2726_ VPWR VGND net1131 sg13g2_dlygate4sd3_1
Xhold363 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[5\] VPWR VGND net1120
+ sg13g2_dlygate4sd3_1
Xhold396 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[5\] VPWR VGND net1153
+ sg13g2_dlygate4sd3_1
X_6209_ _2823_ net508 net1049 VPWR VGND sg13g2_xnor2_1
XFILLER_19_919 VPWR VGND sg13g2_decap_8
XFILLER_45_248 VPWR VGND sg13g2_fill_2
XFILLER_27_974 VPWR VGND sg13g2_decap_8
XFILLER_10_852 VPWR VGND sg13g2_decap_8
XFILLER_6_867 VPWR VGND sg13g2_decap_8
XFILLER_5_377 VPWR VGND sg13g2_fill_2
XFILLER_1_561 VPWR VGND sg13g2_fill_1
XFILLER_18_996 VPWR VGND sg13g2_decap_8
X_3910_ net443 VPWR _0926_ VGND net863 _0925_ sg13g2_o21ai_1
X_4890_ _1730_ _1724_ _1727_ VPWR VGND sg13g2_nand2_1
X_3841_ net419 net875 _0876_ _0021_ VPWR VGND sg13g2_nor3_1
X_6560_ net162 VGND VPWR _0169_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[10\]
+ clknet_leaf_39_clk sg13g2_dfrbpq_1
X_3772_ _0820_ _0539_ net895 VPWR VGND sg13g2_nand2_1
X_5511_ VGND VPWR net524 net1089 _2238_ _2237_ sg13g2_a21oi_1
X_6491_ net231 VGND VPWR _0100_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[5\]
+ clknet_leaf_43_clk sg13g2_dfrbpq_2
X_5442_ _2181_ net1317 _2180_ VPWR VGND sg13g2_nand2_1
X_5373_ net477 VPWR _2123_ VGND _2117_ _2122_ sg13g2_o21ai_1
X_4324_ net770 net436 _0121_ VPWR VGND sg13g2_nor2_1
XFILLER_47_19 VPWR VGND sg13g2_fill_1
X_4255_ VGND VPWR _1194_ _1198_ _1201_ _1197_ sg13g2_a21oi_1
X_4186_ _1142_ _1136_ _1144_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_933 VPWR VGND sg13g2_fill_1
X_6827_ net598 VGND VPWR net1492 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[7\]
+ clknet_leaf_59_clk sg13g2_dfrbpq_2
XFILLER_24_988 VPWR VGND sg13g2_decap_8
X_6758_ net667 VGND VPWR _0367_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[3\]
+ clknet_leaf_31_clk sg13g2_dfrbpq_1
X_5709_ _2400_ _2405_ _2407_ VPWR VGND sg13g2_and2_1
X_6689_ net750 VGND VPWR _0298_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[10\]
+ clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_3_815 VPWR VGND sg13g2_decap_8
Xhold160 _2924_ VPWR VGND net917 sg13g2_dlygate4sd3_1
Xhold171 _0505_ VPWR VGND net928 sg13g2_dlygate4sd3_1
Xhold182 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[0\].z_sign VPWR VGND
+ net939 sg13g2_dlygate4sd3_1
Xhold193 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[2\] VPWR VGND net950 sg13g2_dlygate4sd3_1
XFILLER_46_502 VPWR VGND sg13g2_fill_1
XFILLER_15_955 VPWR VGND sg13g2_decap_8
XFILLER_27_782 VPWR VGND sg13g2_fill_2
X_6477__245 VPWR VGND net245 sg13g2_tiehi
X_4040_ _1033_ _0937_ _1027_ VPWR VGND sg13g2_nand2_1
X_6484__238 VPWR VGND net238 sg13g2_tiehi
XFILLER_18_760 VPWR VGND sg13g2_fill_2
X_5991_ VGND VPWR _2634_ _2636_ _0409_ _2638_ sg13g2_a21oi_1
X_4942_ _1774_ net1160 _1772_ VPWR VGND sg13g2_xnor2_1
X_6612_ net110 VGND VPWR _0221_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[10\]
+ clknet_leaf_24_clk sg13g2_dfrbpq_2
X_4873_ VGND VPWR _0615_ _1710_ _1716_ net536 sg13g2_a21oi_1
XFILLER_21_947 VPWR VGND sg13g2_decap_8
XFILLER_32_251 VPWR VGND sg13g2_fill_1
X_3824_ _0864_ _0862_ _0863_ VPWR VGND sg13g2_xnor2_1
X_6543_ net179 VGND VPWR _0152_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[6\]
+ clknet_leaf_37_clk sg13g2_dfrbpq_2
X_3755_ _0808_ _0797_ _0786_ VPWR VGND sg13g2_nand2b_1
X_6474_ net248 VGND VPWR _0083_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[0\]
+ clknet_leaf_37_clk sg13g2_dfrbpq_2
X_3686_ _0739_ _0738_ _0725_ VPWR VGND sg13g2_nand2b_1
X_5425_ _2166_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[7\] _2165_
+ VPWR VGND sg13g2_xnor2_1
X_5356_ net478 VPWR _2108_ VGND _2103_ _2107_ sg13g2_o21ai_1
XFILLER_0_829 VPWR VGND sg13g2_decap_8
X_4307_ _1246_ net1527 net381 VPWR VGND sg13g2_xnor2_1
X_5287_ net1144 net528 _2050_ VPWR VGND sg13g2_xor2_1
X_4238_ _1187_ net962 net991 VPWR VGND sg13g2_nand2_1
X_4169_ net1356 _1128_ _0097_ VPWR VGND sg13g2_nor2b_1
XFILLER_12_914 VPWR VGND sg13g2_decap_8
XFILLER_11_413 VPWR VGND sg13g2_fill_1
XFILLER_23_251 VPWR VGND sg13g2_fill_1
XFILLER_3_601 VPWR VGND sg13g2_fill_1
XFILLER_3_689 VPWR VGND sg13g2_decap_8
XFILLER_2_144 VPWR VGND sg13g2_fill_2
X_6659__63 VPWR VGND net63 sg13g2_tiehi
Xfanout492 net494 net492 VPWR VGND sg13g2_buf_8
Xfanout481 net482 net481 VPWR VGND sg13g2_buf_8
Xfanout470 net471 net470 VPWR VGND sg13g2_buf_1
XFILLER_0_47 VPWR VGND sg13g2_fill_2
XFILLER_31_1013 VPWR VGND sg13g2_decap_8
X_3540_ VPWR _0610_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[7\] VGND
+ sg13g2_inv_1
XFILLER_7_995 VPWR VGND sg13g2_decap_8
X_3471_ VPWR _0541_ u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[7\] VGND sg13g2_inv_1
X_5210_ _1983_ _1987_ _1988_ VPWR VGND sg13g2_nor2_1
X_6190_ VGND VPWR _0624_ _2795_ _2809_ net510 sg13g2_a21oi_1
X_5141_ _1930_ net493 _1929_ VPWR VGND sg13g2_nand2b_1
X_5072_ net464 VPWR _1882_ VGND _1880_ _1881_ sg13g2_o21ai_1
X_4023_ _1019_ _1018_ _1017_ VPWR VGND sg13g2_nand2b_1
X_5974_ net459 VPWR _2630_ VGND _2628_ _2629_ sg13g2_o21ai_1
X_4925_ net388 net1341 _1760_ VPWR VGND sg13g2_xor2_1
X_4856_ _1702_ net998 net1044 VPWR VGND sg13g2_nand2_1
X_3807_ VGND VPWR net552 _0850_ _0013_ net907 sg13g2_a21oi_1
X_4787_ _1641_ VPWR _1644_ VGND _1637_ _1642_ sg13g2_o21ai_1
X_6526_ net196 VGND VPWR _0135_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[2\]
+ clknet_leaf_39_clk sg13g2_dfrbpq_2
X_3738_ _0791_ net408 _0754_ VPWR VGND sg13g2_xnor2_1
X_3669_ VGND VPWR _0640_ _0703_ _0722_ _0721_ sg13g2_a21oi_1
X_6868__349 VPWR VGND net349 sg13g2_tiehi
X_6457_ net279 VGND VPWR _0066_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[10\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_2
XFILLER_47_1020 VPWR VGND sg13g2_decap_8
X_5408_ net521 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[4\] _2151_
+ VPWR VGND sg13g2_nor2b_1
X_6388_ _0474_ net447 _2891_ _2892_ VPWR VGND sg13g2_and3_1
X_5339_ _2089_ VPWR _2092_ VGND _2086_ _2090_ sg13g2_o21ai_1
XFILLER_0_626 VPWR VGND sg13g2_decap_8
X_6656__66 VPWR VGND net66 sg13g2_tiehi
XFILLER_29_822 VPWR VGND sg13g2_fill_1
XFILLER_18_43 VPWR VGND sg13g2_fill_1
XFILLER_29_899 VPWR VGND sg13g2_fill_1
X_6474__248 VPWR VGND net248 sg13g2_tiehi
X_6851__386 VPWR VGND net570 sg13g2_tiehi
XFILLER_4_965 VPWR VGND sg13g2_decap_8
XFILLER_38_107 VPWR VGND sg13g2_fill_2
XFILLER_38_118 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_58_clk clknet_4_8_0_clk clknet_leaf_58_clk VPWR VGND sg13g2_buf_8
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk VPWR VGND sg13g2_buf_8
X_4710_ _1580_ net1311 _1578_ VPWR VGND sg13g2_xnor2_1
X_5690_ _2388_ net1456 _2390_ VPWR VGND sg13g2_xor2_1
X_4641_ VGND VPWR net537 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[12\]
+ _1522_ _1515_ sg13g2_a21oi_1
X_4572_ VGND VPWR _1459_ _1462_ _1465_ _1464_ sg13g2_a21oi_1
Xhold737 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[3\] VPWR VGND net1494
+ sg13g2_dlygate4sd3_1
XFILLER_7_781 VPWR VGND sg13g2_decap_4
X_3523_ VPWR _0593_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[1\] VGND
+ sg13g2_inv_1
Xhold726 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[6\] VPWR
+ VGND net1483 sg13g2_dlygate4sd3_1
X_6311_ net446 net780 _0485_ VPWR VGND sg13g2_and2_1
Xhold715 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[1\] VPWR
+ VGND net1472 sg13g2_dlygate4sd3_1
Xhold704 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[5\] VPWR VGND net1461
+ sg13g2_dlygate4sd3_1
Xhold748 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[4\] VPWR VGND net1505
+ sg13g2_dlygate4sd3_1
X_6242_ VGND VPWR _2850_ _2849_ _2848_ sg13g2_or2_1
Xhold759 _1680_ VPWR VGND net1516 sg13g2_dlygate4sd3_1
X_6173_ VGND VPWR _0623_ _2780_ _2794_ net507 sg13g2_a21oi_1
X_5124_ _1915_ _1906_ _1913_ VPWR VGND sg13g2_nand2_1
XFILLER_29_107 VPWR VGND sg13g2_fill_2
X_5055_ _1868_ net1219 net395 VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_49_clk clknet_4_11_0_clk clknet_leaf_49_clk VPWR VGND sg13g2_buf_8
X_4006_ _1004_ net954 net376 VPWR VGND sg13g2_nand2_1
X_6653__69 VPWR VGND net69 sg13g2_tiehi
X_6798__443 VPWR VGND net627 sg13g2_tiehi
X_5957_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[11\] net414 _2609_
+ _2615_ VPWR VGND sg13g2_a21o_1
X_4908_ _1746_ net1173 net388 VPWR VGND sg13g2_xnor2_1
X_5888_ net425 net974 _0389_ VPWR VGND sg13g2_nor2_1
X_4839_ _1688_ net1261 _1660_ VPWR VGND sg13g2_nand2_1
X_6509_ net213 VGND VPWR net1529 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[10\]
+ clknet_leaf_44_clk sg13g2_dfrbpq_2
XFILLER_1_924 VPWR VGND sg13g2_decap_8
Xhold20 _0050_ VPWR VGND net777 sg13g2_dlygate4sd3_1
Xhold31 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[9\] VPWR VGND net788
+ sg13g2_dlygate4sd3_1
Xhold42 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[1\] VPWR VGND net799
+ sg13g2_dlygate4sd3_1
Xhold64 u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[8\] VPWR VGND net821 sg13g2_dlygate4sd3_1
Xhold53 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[5\] VPWR VGND net810
+ sg13g2_dlygate4sd3_1
Xhold97 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[15\] VPWR VGND net854
+ sg13g2_dlygate4sd3_1
Xhold86 _0028_ VPWR VGND net843 sg13g2_dlygate4sd3_1
Xhold75 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[10\] VPWR VGND net832
+ sg13g2_dlygate4sd3_1
XFILLER_44_611 VPWR VGND sg13g2_fill_1
XFILLER_44_677 VPWR VGND sg13g2_fill_2
XFILLER_8_589 VPWR VGND sg13g2_fill_2
XFILLER_4_762 VPWR VGND sg13g2_decap_8
XFILLER_6_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_990 VPWR VGND sg13g2_decap_8
X_6860_ net365 VGND VPWR net1042 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[4\]
+ clknet_leaf_64_clk sg13g2_dfrbpq_2
X_5811_ _2483_ VPWR _2489_ VGND net512 _0575_ sg13g2_o21ai_1
XFILLER_16_880 VPWR VGND sg13g2_fill_1
X_6791_ net634 VGND VPWR _0400_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[8\]
+ clknet_leaf_57_clk sg13g2_dfrbpq_2
X_5742_ VGND VPWR net809 _2431_ _2433_ _2430_ sg13g2_a21oi_1
X_5673_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[1\] _2374_
+ _2375_ VPWR VGND sg13g2_and2_1
X_4624_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[8\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[9\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[10\] _1507_ VPWR VGND sg13g2_nor3_1
X_4555_ net1272 net539 _1451_ VPWR VGND sg13g2_xor2_1
Xhold501 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[12\] VPWR VGND net1258
+ sg13g2_dlygate4sd3_1
Xhold545 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[2\] VPWR VGND net1302
+ sg13g2_dlygate4sd3_1
X_3506_ VPWR _0576_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[4\] VGND
+ sg13g2_inv_1
Xhold534 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[11\] VPWR VGND net1291
+ sg13g2_dlygate4sd3_1
X_6910__280 VPWR VGND net280 sg13g2_tiehi
Xhold512 _2065_ VPWR VGND net1269 sg13g2_dlygate4sd3_1
Xhold523 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[2\] VPWR VGND net1280
+ sg13g2_dlygate4sd3_1
Xhold578 _2326_ VPWR VGND net1335 sg13g2_dlygate4sd3_1
Xhold567 _0401_ VPWR VGND net1324 sg13g2_dlygate4sd3_1
Xhold556 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[8\] VPWR VGND net1313
+ sg13g2_dlygate4sd3_1
X_4486_ net543 _1387_ _1394_ VPWR VGND sg13g2_nor2_1
Xhold589 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[7\] VPWR VGND net1346
+ sg13g2_dlygate4sd3_1
X_6225_ net417 net1235 _2836_ VPWR VGND sg13g2_nor2_1
X_6156_ _2772_ VPWR _2779_ VGND net511 _0621_ sg13g2_o21ai_1
X_5107_ VGND VPWR _1890_ _1896_ _1899_ _1895_ sg13g2_a21oi_1
X_6087_ _2719_ net1557 _2720_ VPWR VGND sg13g2_nor2b_1
X_5038_ net470 VPWR _1854_ VGND _1851_ _1852_ sg13g2_o21ai_1
XFILLER_25_187 VPWR VGND sg13g2_fill_2
XFILLER_22_850 VPWR VGND sg13g2_fill_2
Xoutput21 net21 uo_out[4] VPWR VGND sg13g2_buf_1
XFILLER_1_721 VPWR VGND sg13g2_decap_8
XFILLER_1_798 VPWR VGND sg13g2_decap_8
XFILLER_44_463 VPWR VGND sg13g2_fill_1
XFILLER_12_371 VPWR VGND sg13g2_fill_1
XFILLER_9_876 VPWR VGND sg13g2_decap_8
X_6788__453 VPWR VGND net637 sg13g2_tiehi
X_4340_ _1268_ _1271_ _1272_ VPWR VGND sg13g2_and2_1
X_4271_ VGND VPWR _1207_ _1214_ _1216_ net435 sg13g2_a21oi_1
X_6010_ net452 VPWR _2653_ VGND net1046 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[0\]
+ sg13g2_o21ai_1
XFILLER_36_920 VPWR VGND sg13g2_fill_1
X_6912_ net276 VGND VPWR _0507_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[6\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_1
X_6843_ net582 VGND VPWR net969 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[0\]
+ clknet_leaf_64_clk sg13g2_dfrbpq_2
X_6795__446 VPWR VGND net630 sg13g2_tiehi
X_6774_ net651 VGND VPWR net1572 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[7\]
+ clknet_leaf_60_clk sg13g2_dfrbpq_2
X_3986_ _0977_ _0982_ _0984_ _0987_ VGND VPWR _0985_ sg13g2_nor4_2
X_5725_ VGND VPWR _2415_ _2419_ _2421_ net431 sg13g2_a21oi_1
X_5656_ _2359_ net1446 _2360_ VPWR VGND sg13g2_nor2b_1
XFILLER_31_691 VPWR VGND sg13g2_fill_1
X_4607_ net438 net977 _0171_ VPWR VGND sg13g2_nor2_1
X_5587_ VGND VPWR _0595_ _2286_ _2301_ net516 sg13g2_a21oi_1
Xhold320 _0415_ VPWR VGND net1077 sg13g2_dlygate4sd3_1
X_4538_ net385 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[11\] _1438_
+ VPWR VGND sg13g2_xor2_1
Xhold342 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[10\] VPWR VGND net1099
+ sg13g2_dlygate4sd3_1
Xhold353 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[8\] VPWR VGND net1110
+ sg13g2_dlygate4sd3_1
Xhold331 _0167_ VPWR VGND net1088 sg13g2_dlygate4sd3_1
Xhold386 _0197_ VPWR VGND net1143 sg13g2_dlygate4sd3_1
Xhold375 _0426_ VPWR VGND net1132 sg13g2_dlygate4sd3_1
Xhold364 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[9\] VPWR VGND net1121
+ sg13g2_dlygate4sd3_1
X_4469_ _1379_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[0\]
+ net543 VPWR VGND sg13g2_nand2b_1
Xhold397 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[9\] VPWR VGND net1154
+ sg13g2_dlygate4sd3_1
X_6208_ _2822_ _2821_ _0442_ VPWR VGND sg13g2_nor2b_1
X_6139_ VGND VPWR _2757_ _2761_ _2764_ _2760_ sg13g2_a21oi_1
XFILLER_14_603 VPWR VGND sg13g2_fill_1
XFILLER_26_463 VPWR VGND sg13g2_fill_1
X_6917__264 VPWR VGND net264 sg13g2_tiehi
XFILLER_6_846 VPWR VGND sg13g2_decap_8
XFILLER_5_323 VPWR VGND sg13g2_fill_1
XFILLER_49_500 VPWR VGND sg13g2_fill_1
XFILLER_49_555 VPWR VGND sg13g2_fill_2
XFILLER_37_728 VPWR VGND sg13g2_fill_2
XFILLER_18_975 VPWR VGND sg13g2_decap_8
X_3840_ _0876_ net554 net874 net857 VPWR VGND sg13g2_and3_1
X_3771_ VGND VPWR net792 net831 _0008_ _0819_ sg13g2_a21oi_1
XFILLER_20_639 VPWR VGND sg13g2_fill_2
X_5510_ _0329_ net481 _2235_ _2236_ VPWR VGND sg13g2_and3_1
X_6490_ net232 VGND VPWR _0099_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[4\]
+ clknet_leaf_50_clk sg13g2_dfrbpq_2
X_5441_ _2180_ net1570 _2179_ VPWR VGND sg13g2_xnor2_1
X_5372_ _2122_ net1444 _2120_ VPWR VGND sg13g2_xnor2_1
X_4323_ VGND VPWR _1257_ _1258_ _0120_ _1259_ sg13g2_a21oi_1
X_4254_ net1279 _1200_ _0110_ VPWR VGND sg13g2_nor2b_1
X_4185_ _1136_ _1142_ _1143_ VPWR VGND sg13g2_nor2b_1
XFILLER_35_271 VPWR VGND sg13g2_fill_1
X_6826_ net599 VGND VPWR _0435_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[6\]
+ clknet_leaf_59_clk sg13g2_dfrbpq_2
XFILLER_24_967 VPWR VGND sg13g2_decap_8
XFILLER_10_116 VPWR VGND sg13g2_fill_1
X_6757_ net668 VGND VPWR _0366_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[2\]
+ clknet_leaf_29_clk sg13g2_dfrbpq_1
X_5708_ _2400_ _2405_ _2406_ VPWR VGND sg13g2_nor2_1
X_3969_ _0970_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[7\] _0957_
+ VPWR VGND sg13g2_xnor2_1
X_6688_ net751 VGND VPWR net1270 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[9\]
+ clknet_leaf_44_clk sg13g2_dfrbpq_1
X_5639_ VGND VPWR _2341_ _2342_ _2346_ _2343_ sg13g2_a21oi_1
Xhold150 _0849_ VPWR VGND net907 sg13g2_dlygate4sd3_1
Xhold161 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[8\] VPWR VGND
+ net918 sg13g2_dlygate4sd3_1
Xhold183 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[0\] VPWR VGND
+ net940 sg13g2_dlygate4sd3_1
Xhold194 _0877_ VPWR VGND net951 sg13g2_dlygate4sd3_1
Xhold172 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[5\] VPWR VGND net929 sg13g2_dlygate4sd3_1
X_6878__329 VPWR VGND net329 sg13g2_tiehi
XFILLER_15_934 VPWR VGND sg13g2_decap_8
X_6778__463 VPWR VGND net647 sg13g2_tiehi
XFILLER_18_1017 VPWR VGND sg13g2_decap_8
XFILLER_18_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_621 VPWR VGND sg13g2_fill_2
XFILLER_6_632 VPWR VGND sg13g2_fill_2
XFILLER_5_164 VPWR VGND sg13g2_fill_2
X_6785__456 VPWR VGND net640 sg13g2_tiehi
XFILLER_2_893 VPWR VGND sg13g2_decap_8
X_5990_ _2638_ net460 _2637_ VPWR VGND sg13g2_nand2_1
X_4941_ _1773_ net1160 _1772_ VPWR VGND sg13g2_nand2_1
X_4872_ _1714_ VPWR _1715_ VGND _0616_ _1711_ sg13g2_o21ai_1
X_6611_ net111 VGND VPWR net1174 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[9\]
+ clknet_leaf_25_clk sg13g2_dfrbpq_2
X_6792__449 VPWR VGND net633 sg13g2_tiehi
XFILLER_21_926 VPWR VGND sg13g2_decap_8
X_3823_ _0686_ VPWR _0863_ VGND net404 _0755_ sg13g2_o21ai_1
XFILLER_20_425 VPWR VGND sg13g2_fill_1
X_6542_ net180 VGND VPWR _0151_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[5\]
+ clknet_leaf_37_clk sg13g2_dfrbpq_2
XFILLER_9_470 VPWR VGND sg13g2_fill_2
X_3754_ VPWR _0807_ _0806_ VGND sg13g2_inv_1
X_6473_ net249 VGND VPWR _0082_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp\[11\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
X_3685_ _0639_ _0724_ _0637_ _0738_ VPWR VGND sg13g2_nand3_1
X_5424_ VGND VPWR _0558_ _2157_ _2165_ net521 sg13g2_a21oi_1
X_5355_ _2107_ net1417 _2105_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_808 VPWR VGND sg13g2_decap_8
X_4306_ VGND VPWR _1243_ _1244_ _0117_ _1245_ sg13g2_a21oi_1
X_5286_ _2049_ net415 net1144 VPWR VGND sg13g2_nand2_1
X_4237_ VGND VPWR _1184_ _1185_ _0107_ _1186_ sg13g2_a21oi_1
X_4168_ VGND VPWR _1122_ _1126_ _1128_ net439 sg13g2_a21oi_1
X_4099_ net419 _1073_ _0081_ VPWR VGND sg13g2_nor2_1
X_6809_ net616 VGND VPWR net1297 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[4\]
+ clknet_leaf_63_clk sg13g2_dfrbpq_2
XFILLER_48_63 VPWR VGND sg13g2_decap_8
Xfanout493 net494 net493 VPWR VGND sg13g2_buf_1
Xfanout460 net461 net460 VPWR VGND sg13g2_buf_1
Xfanout471 net472 net471 VPWR VGND sg13g2_buf_8
Xfanout482 net490 net482 VPWR VGND sg13g2_buf_1
XFILLER_47_878 VPWR VGND sg13g2_fill_1
XFILLER_46_399 VPWR VGND sg13g2_fill_1
XFILLER_34_528 VPWR VGND sg13g2_decap_4
XFILLER_7_974 VPWR VGND sg13g2_decap_8
X_6490__232 VPWR VGND net232 sg13g2_tiehi
X_3470_ VPWR _0540_ u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[8\] VGND sg13g2_inv_1
XFILLER_43_4 VPWR VGND sg13g2_fill_1
X_5140_ _1926_ _1928_ _1929_ VPWR VGND sg13g2_nor2_1
X_5071_ _1881_ net1197 net396 VPWR VGND sg13g2_xnor2_1
XFILLER_2_690 VPWR VGND sg13g2_decap_8
X_4022_ _1018_ net961 net549 VPWR VGND sg13g2_nand2_1
X_6599__123 VPWR VGND net123 sg13g2_tiehi
X_5973_ _2622_ net1323 _2629_ VPWR VGND sg13g2_xor2_1
XFILLER_37_399 VPWR VGND sg13g2_fill_1
X_4924_ net1565 _1759_ _0221_ VPWR VGND sg13g2_nor2_1
X_4855_ VGND VPWR _1699_ _1700_ _0210_ _1701_ sg13g2_a21oi_1
X_4786_ VGND VPWR _1637_ _1642_ _0199_ _1643_ sg13g2_a21oi_1
X_3806_ _0850_ _0747_ _0768_ VPWR VGND sg13g2_xnor2_1
X_6525_ net197 VGND VPWR net1098 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[1\]
+ clknet_leaf_38_clk sg13g2_dfrbpq_1
X_3737_ _0790_ net408 _0754_ VPWR VGND sg13g2_nand2_1
X_3668_ _0719_ _0720_ _0721_ VPWR VGND sg13g2_nor2_1
X_6456_ net281 VGND VPWR net1013 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[9\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_2
X_5407_ net439 net1055 _0313_ VPWR VGND sg13g2_nor2_1
X_6387_ VGND VPWR _2857_ _2882_ _0469_ _2886_ sg13g2_a21oi_1
X_3599_ _0652_ _0636_ _0651_ VPWR VGND sg13g2_nand2_1
X_5338_ VGND VPWR _2086_ net1256 _0303_ _2091_ sg13g2_a21oi_1
X_6768__473 VPWR VGND net657 sg13g2_tiehi
X_5269_ net804 net435 _0290_ VPWR VGND sg13g2_nor2_1
X_6699__556 VPWR VGND net740 sg13g2_tiehi
XFILLER_24_550 VPWR VGND sg13g2_fill_1
X_6775__466 VPWR VGND net650 sg13g2_tiehi
XFILLER_34_87 VPWR VGND sg13g2_fill_2
XFILLER_4_944 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_fill_2
X_6450__293 VPWR VGND net293 sg13g2_tiehi
X_6782__459 VPWR VGND net643 sg13g2_tiehi
XFILLER_46_163 VPWR VGND sg13g2_fill_1
X_4640_ VGND VPWR _1513_ _1519_ _0175_ _1521_ sg13g2_a21oi_1
XFILLER_7_760 VPWR VGND sg13g2_decap_8
X_6310_ net446 net778 _0484_ VPWR VGND sg13g2_and2_1
X_4571_ net1153 net539 _1464_ VPWR VGND sg13g2_xor2_1
Xhold705 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[7\] VPWR VGND net1462
+ sg13g2_dlygate4sd3_1
X_3522_ _0592_ net519 VPWR VGND sg13g2_inv_2
Xhold727 _2220_ VPWR VGND net1484 sg13g2_dlygate4sd3_1
Xhold716 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[5\] VPWR VGND net1473
+ sg13g2_dlygate4sd3_1
Xhold738 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[6\] VPWR VGND net1495
+ sg13g2_dlygate4sd3_1
X_6241_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[9\] net510 _2849_
+ VPWR VGND sg13g2_xor2_1
Xhold749 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[6\] VPWR VGND net1506
+ sg13g2_dlygate4sd3_1
X_6172_ _2790_ _2786_ _2789_ _2793_ VPWR VGND sg13g2_a21o_1
X_5123_ _1914_ _1912_ _1906_ VPWR VGND sg13g2_nand2b_1
XFILLER_34_0 VPWR VGND sg13g2_fill_2
X_5054_ VGND VPWR u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[7\] _1843_
+ _1867_ _1866_ sg13g2_a21oi_1
X_4005_ _0999_ VPWR _0058_ VGND net372 _1003_ sg13g2_o21ai_1
X_5956_ _2614_ _2613_ _0398_ VPWR VGND sg13g2_nor2b_1
X_4907_ _1745_ net1173 net388 VPWR VGND sg13g2_nand2_1
X_5887_ _2555_ net973 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[2\]
+ VPWR VGND sg13g2_xnor2_1
X_4838_ VGND VPWR _1684_ _1686_ _0207_ _1687_ sg13g2_a21oi_1
X_6397__383 VPWR VGND net567 sg13g2_tiehi
X_4769_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[2\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[1\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[3\] _1629_ VPWR VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[0\]
+ sg13g2_nand4_1
X_6508_ net214 VGND VPWR net1513 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[9\]
+ clknet_leaf_41_clk sg13g2_dfrbpq_2
X_6439_ net308 VGND VPWR _0048_ u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[5\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_1_903 VPWR VGND sg13g2_decap_8
Xhold21 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[7\] VPWR VGND net778
+ sg13g2_dlygate4sd3_1
Xhold10 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[1\] VPWR VGND net767
+ sg13g2_dlygate4sd3_1
Xhold32 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[10\] VPWR VGND net789
+ sg13g2_dlygate4sd3_1
Xhold65 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.x_start\[0\] VPWR VGND
+ net822 sg13g2_dlygate4sd3_1
Xhold54 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[10\] VPWR VGND net811
+ sg13g2_dlygate4sd3_1
XFILLER_29_65 VPWR VGND sg13g2_fill_2
Xhold43 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[0\] VPWR VGND net800
+ sg13g2_dlygate4sd3_1
Xhold98 _0516_ VPWR VGND net855 sg13g2_dlygate4sd3_1
XFILLER_21_1024 VPWR VGND sg13g2_decap_4
Xhold87 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[5\] VPWR VGND net844
+ sg13g2_dlygate4sd3_1
Xhold76 _0170_ VPWR VGND net833 sg13g2_dlygate4sd3_1
X_6652__70 VPWR VGND net70 sg13g2_tiehi
X_6480__242 VPWR VGND net242 sg13g2_tiehi
XFILLER_43_155 VPWR VGND sg13g2_fill_2
X_6406__368 VPWR VGND net368 sg13g2_tiehi
XFILLER_8_502 VPWR VGND sg13g2_fill_1
XFILLER_12_586 VPWR VGND sg13g2_fill_1
XFILLER_4_741 VPWR VGND sg13g2_decap_8
X_6589__133 VPWR VGND net133 sg13g2_tiehi
XFILLER_6_1007 VPWR VGND sg13g2_decap_8
X_5810_ net1475 VPWR _2488_ VGND _2482_ _2486_ sg13g2_o21ai_1
XFILLER_16_870 VPWR VGND sg13g2_fill_1
X_6790_ net635 VGND VPWR _0399_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[7\]
+ clknet_leaf_58_clk sg13g2_dfrbpq_2
XFILLER_34_155 VPWR VGND sg13g2_fill_1
X_6596__126 VPWR VGND net126 sg13g2_tiehi
X_5741_ VGND VPWR net809 _2431_ _0365_ _2432_ sg13g2_a21oi_1
X_6758__483 VPWR VGND net667 sg13g2_tiehi
X_5672_ _2372_ net1401 _2374_ VPWR VGND sg13g2_xor2_1
XFILLER_31_895 VPWR VGND sg13g2_fill_2
X_4623_ VGND VPWR _1498_ _1503_ _1506_ _1502_ sg13g2_a21oi_1
X_4554_ _1450_ _1449_ _0160_ VPWR VGND sg13g2_nor2b_1
Xhold502 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[7\] VPWR VGND net1259
+ sg13g2_dlygate4sd3_1
X_3505_ VPWR _0575_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[2\]
+ VGND sg13g2_inv_1
Xhold524 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[11\] VPWR
+ VGND net1281 sg13g2_dlygate4sd3_1
Xhold535 _0273_ VPWR VGND net1292 sg13g2_dlygate4sd3_1
Xhold513 _0297_ VPWR VGND net1270 sg13g2_dlygate4sd3_1
Xhold546 _0340_ VPWR VGND net1303 sg13g2_dlygate4sd3_1
Xhold579 _0346_ VPWR VGND net1336 sg13g2_dlygate4sd3_1
Xhold557 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[6\] VPWR
+ VGND net1314 sg13g2_dlygate4sd3_1
X_6224_ _2831_ _2834_ _2835_ VPWR VGND sg13g2_and2_1
Xhold568 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[8\] VPWR VGND net1325
+ sg13g2_dlygate4sd3_1
X_6689__566 VPWR VGND net750 sg13g2_tiehi
X_4485_ VGND VPWR _1384_ _1390_ _1393_ _1389_ sg13g2_a21oi_1
X_6155_ _2776_ _2770_ _2774_ _2778_ VPWR VGND sg13g2_a21o_1
X_6086_ _2719_ _0625_ _2718_ VPWR VGND sg13g2_xnor2_1
X_5106_ net1394 _1898_ _0264_ VPWR VGND sg13g2_nor2b_1
X_6765__476 VPWR VGND net660 sg13g2_tiehi
X_5037_ VPWR _1853_ _1852_ VGND sg13g2_inv_1
XFILLER_26_623 VPWR VGND sg13g2_decap_8
XFILLER_26_645 VPWR VGND sg13g2_fill_1
XFILLER_41_604 VPWR VGND sg13g2_fill_2
X_6696__559 VPWR VGND net743 sg13g2_tiehi
XFILLER_41_637 VPWR VGND sg13g2_fill_1
X_5939_ _2600_ _0577_ _2598_ VPWR VGND sg13g2_xnor2_1
X_6772__469 VPWR VGND net653 sg13g2_tiehi
XFILLER_22_884 VPWR VGND sg13g2_fill_2
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk VPWR VGND sg13g2_buf_8
XFILLER_1_700 VPWR VGND sg13g2_decap_8
Xoutput22 net22 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_777 VPWR VGND sg13g2_decap_8
XFILLER_44_453 VPWR VGND sg13g2_fill_2
XFILLER_13_851 VPWR VGND sg13g2_fill_2
X_6857__371 VPWR VGND net371 sg13g2_tiehi
XFILLER_13_895 VPWR VGND sg13g2_decap_8
XFILLER_40_670 VPWR VGND sg13g2_fill_2
XFILLER_9_855 VPWR VGND sg13g2_decap_8
X_4270_ _1207_ _1214_ _1215_ VPWR VGND sg13g2_nor2_1
XFILLER_11_2 VPWR VGND sg13g2_fill_1
XFILLER_48_770 VPWR VGND sg13g2_fill_1
X_6911_ net278 VGND VPWR net845 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[5\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_2
X_6842_ net583 VGND VPWR _0451_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].z_sign
+ clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_35_475 VPWR VGND sg13g2_fill_1
XFILLER_36_987 VPWR VGND sg13g2_fill_2
X_6773_ net652 VGND VPWR net1308 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[6\]
+ clknet_leaf_60_clk sg13g2_dfrbpq_2
X_3985_ _0977_ _0982_ _0984_ _0986_ VGND VPWR _0985_ sg13g2_nor4_2
X_5724_ _2415_ _2419_ _2420_ VPWR VGND sg13g2_nor2_1
X_5655_ _2359_ _0596_ _2358_ VPWR VGND sg13g2_xnor2_1
X_4606_ _1492_ net976 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[8\]
+ VPWR VGND sg13g2_xnor2_1
Xhold310 _0010_ VPWR VGND net1067 sg13g2_dlygate4sd3_1
X_5586_ _2297_ VPWR _2300_ VGND _2293_ _2298_ sg13g2_o21ai_1
X_4537_ net438 _1436_ _1437_ _0156_ VPWR VGND sg13g2_nor3_1
Xhold343 _2856_ VPWR VGND net1100 sg13g2_dlygate4sd3_1
Xhold321 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[7\] VPWR VGND net1078
+ sg13g2_dlygate4sd3_1
Xhold332 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[3\] VPWR VGND net1089
+ sg13g2_dlygate4sd3_1
X_4468_ net986 _1377_ _0146_ VPWR VGND sg13g2_nor2b_1
Xhold387 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[6\] VPWR VGND net1144
+ sg13g2_dlygate4sd3_1
Xhold365 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[6\] VPWR VGND net1122
+ sg13g2_dlygate4sd3_1
Xhold376 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[7\] VPWR VGND net1133
+ sg13g2_dlygate4sd3_1
Xhold354 _0129_ VPWR VGND net1111 sg13g2_dlygate4sd3_1
Xhold398 _0411_ VPWR VGND net1155 sg13g2_dlygate4sd3_1
X_6207_ net466 VPWR _2822_ VGND net759 _2820_ sg13g2_o21ai_1
X_6138_ _2762_ _2763_ _0431_ VPWR VGND sg13g2_nor2b_1
X_4399_ _1317_ _1311_ _1315_ _1320_ VPWR VGND sg13g2_a21o_1
X_6069_ _2705_ net452 _2704_ VPWR VGND sg13g2_nand2_1
XFILLER_14_637 VPWR VGND sg13g2_fill_2
X_6579__143 VPWR VGND net143 sg13g2_tiehi
XFILLER_13_147 VPWR VGND sg13g2_fill_2
XFILLER_6_825 VPWR VGND sg13g2_decap_8
XFILLER_10_887 VPWR VGND sg13g2_decap_8
X_6586__136 VPWR VGND net136 sg13g2_tiehi
XFILLER_1_541 VPWR VGND sg13g2_fill_2
X_6748__493 VPWR VGND net677 sg13g2_tiehi
XFILLER_18_954 VPWR VGND sg13g2_decap_8
XFILLER_33_968 VPWR VGND sg13g2_fill_1
X_3770_ net441 VPWR _0819_ VGND net792 net831 sg13g2_o21ai_1
XFILLER_32_478 VPWR VGND sg13g2_fill_2
X_6593__129 VPWR VGND net129 sg13g2_tiehi
X_6755__486 VPWR VGND net670 sg13g2_tiehi
X_5440_ VGND VPWR _0560_ _2172_ _2179_ net521 sg13g2_a21oi_1
X_5371_ _2121_ net1444 _2120_ VPWR VGND sg13g2_nand2_1
XFILLER_5_891 VPWR VGND sg13g2_decap_8
X_4322_ net497 VPWR _1259_ VGND _1257_ _1258_ sg13g2_o21ai_1
X_4253_ VGND VPWR _1194_ _1198_ _1200_ net429 sg13g2_a21oi_1
X_6686__569 VPWR VGND net753 sg13g2_tiehi
X_4184_ _1142_ _1141_ _1140_ VPWR VGND sg13g2_nand2b_1
X_6762__479 VPWR VGND net663 sg13g2_tiehi
XFILLER_24_946 VPWR VGND sg13g2_decap_8
X_6825_ net600 VGND VPWR _0434_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[5\]
+ clknet_leaf_59_clk sg13g2_dfrbpq_1
X_3968_ _0969_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[11\] _0968_
+ VPWR VGND sg13g2_xnor2_1
X_6756_ net669 VGND VPWR _0365_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[1\]
+ clknet_leaf_31_clk sg13g2_dfrbpq_1
X_5707_ VPWR _2405_ _2404_ VGND sg13g2_inv_1
X_3899_ net420 net942 _0918_ _0037_ VPWR VGND sg13g2_nor3_1
X_6687_ net752 VGND VPWR _0296_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[8\]
+ clknet_leaf_43_clk sg13g2_dfrbpq_1
X_5638_ VGND VPWR _2341_ _2344_ _0349_ _2345_ sg13g2_a21oi_1
X_5569_ VGND VPWR _0594_ _2278_ _2285_ net515 sg13g2_a21oi_1
Xhold140 _0009_ VPWR VGND net897 sg13g2_dlygate4sd3_1
Xhold151 _0013_ VPWR VGND net908 sg13g2_dlygate4sd3_1
Xhold162 u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[2\] VPWR VGND net919 sg13g2_dlygate4sd3_1
Xhold173 _0004_ VPWR VGND net930 sg13g2_dlygate4sd3_1
Xhold184 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[6\] VPWR VGND net941 sg13g2_dlygate4sd3_1
Xhold195 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[6\] VPWR VGND
+ net952 sg13g2_dlygate4sd3_1
XFILLER_15_913 VPWR VGND sg13g2_decap_8
XFILLER_30_949 VPWR VGND sg13g2_fill_1
XFILLER_2_872 VPWR VGND sg13g2_decap_8
XFILLER_49_397 VPWR VGND sg13g2_fill_2
X_4940_ _1772_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[11\] _1771_
+ VPWR VGND sg13g2_xnor2_1
X_4871_ _0213_ net484 _1713_ _1714_ VPWR VGND sg13g2_and3_1
XFILLER_33_765 VPWR VGND sg13g2_fill_1
X_6610_ net112 VGND VPWR _0219_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[8\]
+ clknet_leaf_24_clk sg13g2_dfrbpq_1
X_3822_ VGND VPWR _0862_ _0861_ _0860_ sg13g2_or2_1
X_6541_ net181 VGND VPWR _0150_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[4\]
+ clknet_leaf_35_clk sg13g2_dfrbpq_1
XFILLER_14_990 VPWR VGND sg13g2_decap_8
X_3753_ _0806_ _0800_ _0804_ VPWR VGND sg13g2_xnor2_1
X_6472_ net251 VGND VPWR _0081_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[11\]
+ clknet_leaf_0_clk sg13g2_dfrbpq_2
X_3684_ _0733_ _0736_ _0737_ VPWR VGND sg13g2_nor2_1
X_5423_ VGND VPWR _2156_ _2161_ _2164_ _2160_ sg13g2_a21oi_1
X_5354_ _2106_ net1417 _2105_ VPWR VGND sg13g2_nand2_1
X_6668__54 VPWR VGND net54 sg13g2_tiehi
X_4305_ net501 VPWR _1245_ VGND _1243_ _1244_ sg13g2_o21ai_1
X_5285_ _2044_ _2047_ _2048_ VPWR VGND sg13g2_and2_1
X_6569__153 VPWR VGND net153 sg13g2_tiehi
X_4236_ net496 VPWR _1186_ VGND _1184_ _1185_ sg13g2_o21ai_1
X_4167_ _1122_ _1126_ _1127_ VPWR VGND sg13g2_nor2_1
X_6907__286 VPWR VGND net286 sg13g2_tiehi
XFILLER_28_548 VPWR VGND sg13g2_fill_1
XFILLER_43_507 VPWR VGND sg13g2_fill_1
X_4098_ _1072_ net878 _1073_ VPWR VGND sg13g2_xor2_1
XFILLER_43_529 VPWR VGND sg13g2_fill_2
X_6808_ net617 VGND VPWR net1340 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[3\]
+ clknet_leaf_62_clk sg13g2_dfrbpq_2
XFILLER_24_787 VPWR VGND sg13g2_fill_1
XFILLER_8_909 VPWR VGND sg13g2_decap_8
XFILLER_12_949 VPWR VGND sg13g2_decap_8
X_6576__146 VPWR VGND net146 sg13g2_tiehi
X_6739_ net686 VGND VPWR net1469 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[10\]
+ clknet_leaf_57_clk sg13g2_dfrbpq_2
XFILLER_20_982 VPWR VGND sg13g2_decap_8
XFILLER_2_102 VPWR VGND sg13g2_fill_1
XFILLER_48_42 VPWR VGND sg13g2_decap_8
Xfanout450 net451 net450 VPWR VGND sg13g2_buf_8
X_6583__139 VPWR VGND net139 sg13g2_tiehi
Xfanout461 net473 net461 VPWR VGND sg13g2_buf_2
Xfanout472 net473 net472 VPWR VGND sg13g2_buf_8
Xfanout483 net485 net483 VPWR VGND sg13g2_buf_8
X_6745__496 VPWR VGND net680 sg13g2_tiehi
Xfanout494 net495 net494 VPWR VGND sg13g2_buf_1
XFILLER_15_787 VPWR VGND sg13g2_fill_1
XFILLER_15_798 VPWR VGND sg13g2_fill_2
X_6791__450 VPWR VGND net634 sg13g2_tiehi
XFILLER_7_953 VPWR VGND sg13g2_decap_8
XFILLER_11_982 VPWR VGND sg13g2_decap_8
X_6752__489 VPWR VGND net673 sg13g2_tiehi
X_6416__348 VPWR VGND net348 sg13g2_tiehi
XFILLER_9_1016 VPWR VGND sg13g2_decap_8
XFILLER_9_1027 VPWR VGND sg13g2_fill_2
XFILLER_36_4 VPWR VGND sg13g2_fill_2
X_5070_ _1878_ VPWR _1880_ VGND _0544_ net396 sg13g2_o21ai_1
X_6665__57 VPWR VGND net57 sg13g2_tiehi
X_4021_ net961 net549 _1017_ VPWR VGND sg13g2_nor2_1
X_5972_ VGND VPWR _2620_ _2623_ _2628_ _2627_ sg13g2_a21oi_1
XFILLER_25_518 VPWR VGND sg13g2_fill_2
X_4923_ _1759_ net483 _1758_ VPWR VGND sg13g2_nand2_1
XFILLER_18_581 VPWR VGND sg13g2_decap_8
XFILLER_33_551 VPWR VGND sg13g2_fill_1
XFILLER_33_562 VPWR VGND sg13g2_fill_1
X_4854_ net483 VPWR _1701_ VGND _1699_ _1700_ sg13g2_o21ai_1
X_4785_ net485 VPWR _1643_ VGND _1637_ _1642_ sg13g2_o21ai_1
X_3805_ net552 net906 _0849_ VPWR VGND sg13g2_nor2_1
X_6524_ net198 VGND VPWR _0133_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[0\]
+ clknet_leaf_38_clk sg13g2_dfrbpq_1
X_3736_ _0777_ VPWR _0789_ VGND _0776_ _0779_ sg13g2_o21ai_1
X_3667_ _0720_ _0640_ _0703_ VPWR VGND sg13g2_xnor2_1
X_6455_ net283 VGND VPWR _0064_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[8\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_2
X_5406_ _2150_ net1054 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[4\]
+ VPWR VGND sg13g2_xnor2_1
X_6386_ VGND VPWR net402 _2882_ _0468_ _2886_ sg13g2_a21oi_1
X_3598_ _0649_ _0650_ _0651_ VPWR VGND _0648_ sg13g2_nand3b_1
X_5337_ net477 VPWR _2091_ VGND _2086_ _2090_ sg13g2_o21ai_1
X_5268_ net489 net830 _0289_ VPWR VGND sg13g2_and2_1
X_4219_ VGND VPWR _1169_ _1170_ _0104_ _1171_ sg13g2_a21oi_1
X_5199_ _1978_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[8\] _1977_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_43_359 VPWR VGND sg13g2_fill_1
XFILLER_7_205 VPWR VGND sg13g2_fill_1
XFILLER_4_923 VPWR VGND sg13g2_decap_8
X_6559__163 VPWR VGND net163 sg13g2_tiehi
X_4570_ VGND VPWR _1460_ _1461_ _0163_ _1463_ sg13g2_a21oi_1
X_3521_ VPWR _0591_ net1115 VGND sg13g2_inv_1
Xhold717 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[2\] VPWR VGND net1474
+ sg13g2_dlygate4sd3_1
Xhold728 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[3\] VPWR VGND net1485
+ sg13g2_dlygate4sd3_1
Xhold706 _1237_ VPWR VGND net1463 sg13g2_dlygate4sd3_1
Xhold739 _1599_ VPWR VGND net1496 sg13g2_dlygate4sd3_1
X_6240_ VGND VPWR net508 net1071 _2848_ _2846_ sg13g2_a21oi_1
X_6171_ _2791_ _2792_ _0435_ VPWR VGND sg13g2_nor2b_1
X_6867__351 VPWR VGND net351 sg13g2_tiehi
X_5122_ VPWR _1913_ _1912_ VGND sg13g2_inv_1
X_5053_ _1866_ _1855_ _1857_ VPWR VGND sg13g2_nand2_1
X_6566__156 VPWR VGND net156 sg13g2_tiehi
X_4004_ _1003_ _1002_ _1001_ VPWR VGND sg13g2_nand2b_1
X_5955_ net459 VPWR _2614_ VGND _2608_ _2612_ sg13g2_o21ai_1
X_4906_ _1741_ _1743_ _1744_ VPWR VGND sg13g2_nor2_1
X_5886_ net973 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[2\] _2554_
+ VPWR VGND sg13g2_nor2b_1
X_4837_ net471 VPWR _1687_ VGND _1684_ _1686_ sg13g2_o21ai_1
X_4768_ VGND VPWR _1626_ _1627_ _0196_ _1628_ sg13g2_a21oi_1
XFILLER_5_709 VPWR VGND sg13g2_decap_8
X_6573__149 VPWR VGND net149 sg13g2_tiehi
X_3719_ VGND VPWR _0771_ _0772_ _0770_ _0744_ sg13g2_a21oi_2
X_6507_ net215 VGND VPWR _0116_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[8\]
+ clknet_leaf_44_clk sg13g2_dfrbpq_2
X_4699_ net537 _1549_ _1570_ VPWR VGND sg13g2_nor2_1
X_6438_ net309 VGND VPWR _0047_ u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[4\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_20_79 VPWR VGND sg13g2_fill_2
XFILLER_1_959 VPWR VGND sg13g2_decap_8
X_6369_ _2921_ _2922_ _0515_ VPWR VGND sg13g2_nor2_1
Xhold22 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[2\] VPWR VGND net779
+ sg13g2_dlygate4sd3_1
Xhold11 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[1\] VPWR VGND net768
+ sg13g2_dlygate4sd3_1
Xhold33 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[2\] VPWR VGND net790
+ sg13g2_dlygate4sd3_1
X_6781__460 VPWR VGND net644 sg13g2_tiehi
Xhold55 _0337_ VPWR VGND net812 sg13g2_dlygate4sd3_1
Xhold44 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[5\] VPWR VGND net801
+ sg13g2_dlygate4sd3_1
Xhold66 _0003_ VPWR VGND net823 sg13g2_dlygate4sd3_1
Xhold99 u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[6\] VPWR VGND net856 sg13g2_dlygate4sd3_1
XFILLER_21_1003 VPWR VGND sg13g2_decap_8
Xhold88 _0506_ VPWR VGND net845 sg13g2_dlygate4sd3_1
Xhold77 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[2\] VPWR VGND net834
+ sg13g2_dlygate4sd3_1
XFILLER_43_134 VPWR VGND sg13g2_fill_1
XFILLER_43_101 VPWR VGND sg13g2_fill_1
X_6742__499 VPWR VGND net683 sg13g2_tiehi
XFILLER_12_510 VPWR VGND sg13g2_fill_1
XFILLER_24_381 VPWR VGND sg13g2_fill_2
XFILLER_4_720 VPWR VGND sg13g2_decap_8
XFILLER_4_797 VPWR VGND sg13g2_decap_8
XFILLER_39_429 VPWR VGND sg13g2_fill_2
XFILLER_34_145 VPWR VGND sg13g2_fill_1
XFILLER_16_893 VPWR VGND sg13g2_decap_8
X_5740_ net468 VPWR _2432_ VGND net809 _2431_ sg13g2_o21ai_1
X_5671_ _2373_ _2372_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[7\]
+ VPWR VGND sg13g2_nand2b_1
X_4622_ _1504_ _1505_ _0173_ VPWR VGND sg13g2_nor2b_1
X_4553_ net502 VPWR _1450_ VGND net760 _1448_ sg13g2_o21ai_1
Xhold503 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[9\] VPWR VGND net1260
+ sg13g2_dlygate4sd3_1
Xhold536 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[5\] VPWR VGND net1293
+ sg13g2_dlygate4sd3_1
X_3504_ VPWR _0574_ net1427 VGND sg13g2_inv_1
Xhold525 _2817_ VPWR VGND net1282 sg13g2_dlygate4sd3_1
Xhold514 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[5\] VPWR VGND net1271
+ sg13g2_dlygate4sd3_1
X_4484_ net1225 _1392_ _0148_ VPWR VGND sg13g2_nor2b_1
Xhold547 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[4\]\[1\] VPWR VGND net1304
+ sg13g2_dlygate4sd3_1
Xhold569 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[9\] VPWR VGND net1326
+ sg13g2_dlygate4sd3_1
Xhold558 _2033_ VPWR VGND net1315 sg13g2_dlygate4sd3_1
X_6223_ _0445_ net455 net1330 _2834_ VPWR VGND sg13g2_and3_1
X_6154_ VGND VPWR _2771_ _2775_ _0433_ _2777_ sg13g2_a21oi_1
X_6085_ VGND VPWR net417 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[9\]
+ _2718_ _2712_ sg13g2_a21oi_1
X_5105_ VGND VPWR _1890_ _1896_ _1898_ net430 sg13g2_a21oi_1
X_5036_ _1852_ net1396 net396 VPWR VGND sg13g2_xnor2_1
XFILLER_38_484 VPWR VGND sg13g2_fill_2
X_5938_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[5\] _2598_
+ _2599_ VPWR VGND sg13g2_and2_1
X_5869_ VGND VPWR net413 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[9\]
+ _2540_ _2534_ sg13g2_a21oi_1
Xoutput23 net23 uo_out[7] VPWR VGND sg13g2_buf_1
XFILLER_0_211 VPWR VGND sg13g2_fill_2
XFILLER_1_756 VPWR VGND sg13g2_decap_8
X_6549__173 VPWR VGND net173 sg13g2_tiehi
XFILLER_45_999 VPWR VGND sg13g2_fill_1
XFILLER_17_679 VPWR VGND sg13g2_fill_1
XFILLER_12_395 VPWR VGND sg13g2_fill_2
X_6556__166 VPWR VGND net166 sg13g2_tiehi
X_6563__159 VPWR VGND net159 sg13g2_tiehi
X_6910_ net280 VGND VPWR net928 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[4\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_35_410 VPWR VGND sg13g2_fill_2
X_6841_ net584 VGND VPWR _0450_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[10\]
+ clknet_leaf_9_clk sg13g2_dfrbpq_1
X_6772_ net653 VGND VPWR _0381_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[5\]
+ clknet_leaf_60_clk sg13g2_dfrbpq_1
X_6695__560 VPWR VGND net744 sg13g2_tiehi
X_3984_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[16\] _0983_ _0985_
+ VPWR VGND sg13g2_nor2b_2
X_5723_ VPWR _2419_ _2418_ VGND sg13g2_inv_1
X_5654_ net515 _2357_ _2358_ VPWR VGND sg13g2_nor2_1
X_4605_ net976 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[8\] _1491_
+ VPWR VGND sg13g2_nor2b_1
X_6771__470 VPWR VGND net654 sg13g2_tiehi
X_5585_ VGND VPWR _2293_ _2298_ _0342_ _2299_ sg13g2_a21oi_1
XFILLER_11_1024 VPWR VGND sg13g2_decap_4
Xhold311 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[10\] VPWR VGND net1068
+ sg13g2_dlygate4sd3_1
Xhold300 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[3\] VPWR VGND net1057
+ sg13g2_dlygate4sd3_1
Xhold344 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[0\] VPWR
+ VGND net1101 sg13g2_dlygate4sd3_1
Xhold322 _0371_ VPWR VGND net1079 sg13g2_dlygate4sd3_1
Xhold333 _0330_ VPWR VGND net1090 sg13g2_dlygate4sd3_1
X_4536_ VGND VPWR _1433_ _1434_ _1437_ _1435_ sg13g2_a21oi_1
X_4467_ net486 VPWR _1378_ VGND net985 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[0\]
+ sg13g2_o21ai_1
Xhold366 _0231_ VPWR VGND net1123 sg13g2_dlygate4sd3_1
Xhold355 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[4\] VPWR VGND net1112
+ sg13g2_dlygate4sd3_1
Xhold377 _1474_ VPWR VGND net1134 sg13g2_dlygate4sd3_1
Xhold399 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[7\] VPWR VGND net1156
+ sg13g2_dlygate4sd3_1
X_6206_ _2821_ net759 _2820_ VPWR VGND sg13g2_nand2_1
Xhold388 _0294_ VPWR VGND net1145 sg13g2_dlygate4sd3_1
X_4398_ _1318_ _1319_ _0135_ VPWR VGND sg13g2_nor2b_1
X_6137_ VGND VPWR _2757_ _2761_ _2763_ net422 sg13g2_a21oi_1
X_6068_ _2702_ VPWR _2704_ VGND _2691_ _2695_ sg13g2_o21ai_1
X_5019_ _1838_ net1488 _1836_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_12 VPWR VGND sg13g2_fill_1
XFILLER_26_421 VPWR VGND sg13g2_fill_1
XFILLER_27_988 VPWR VGND sg13g2_decap_8
XFILLER_26_487 VPWR VGND sg13g2_fill_2
XFILLER_41_424 VPWR VGND sg13g2_fill_1
XFILLER_13_159 VPWR VGND sg13g2_fill_2
XFILLER_6_804 VPWR VGND sg13g2_decap_8
XFILLER_10_866 VPWR VGND sg13g2_decap_8
XFILLER_18_933 VPWR VGND sg13g2_decap_8
X_6447__299 VPWR VGND net299 sg13g2_tiehi
X_5370_ _2120_ _0559_ _2119_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_870 VPWR VGND sg13g2_decap_8
X_4321_ _1258_ net1199 net381 VPWR VGND sg13g2_xnor2_1
X_4252_ _1194_ net1278 _1199_ VPWR VGND sg13g2_nor2_1
X_4183_ _1141_ _1139_ net1499 VPWR VGND sg13g2_nand2b_1
X_6426__328 VPWR VGND net328 sg13g2_tiehi
X_6824_ net601 VGND VPWR _0433_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[4\]
+ clknet_leaf_60_clk sg13g2_dfrbpq_2
X_3967_ _0944_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[6\] _0968_
+ VPWR VGND sg13g2_xor2_1
X_6755_ net670 VGND VPWR _0364_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[0\]
+ clknet_leaf_29_clk sg13g2_dfrbpq_2
X_5706_ _2404_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[5\]
+ _2402_ VPWR VGND sg13g2_xnor2_1
X_3898_ _0918_ net941 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[5\] _0915_ VPWR VGND
+ sg13g2_and3_2
Xclkbuf_leaf_30_clk clknet_4_9_0_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
X_6686_ net753 VGND VPWR _0295_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[7\]
+ clknet_leaf_44_clk sg13g2_dfrbpq_1
X_6539__183 VPWR VGND net183 sg13g2_tiehi
X_5637_ net476 VPWR _2345_ VGND _2341_ _2344_ sg13g2_o21ai_1
XFILLER_3_829 VPWR VGND sg13g2_decap_8
X_5568_ _2281_ VPWR _2284_ VGND _2277_ _2282_ sg13g2_o21ai_1
X_4519_ _1423_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[7\] net384
+ VPWR VGND sg13g2_xnor2_1
Xhold130 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[9\] VPWR VGND net887 sg13g2_dlygate4sd3_1
Xhold152 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[3\] VPWR VGND net909 sg13g2_dlygate4sd3_1
Xhold141 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[2\] VPWR VGND net898
+ sg13g2_dlygate4sd3_1
Xhold163 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[2\] VPWR VGND net920 sg13g2_dlygate4sd3_1
Xhold185 _0917_ VPWR VGND net942 sg13g2_dlygate4sd3_1
Xhold174 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[3\] VPWR VGND net931
+ sg13g2_dlygate4sd3_1
X_5499_ VGND VPWR net852 _2227_ _0327_ _2228_ sg13g2_a21oi_1
Xhold196 _0062_ VPWR VGND net953 sg13g2_dlygate4sd3_1
X_6546__176 VPWR VGND net176 sg13g2_tiehi
XFILLER_15_969 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_21_clk clknet_4_5_0_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
X_6592__130 VPWR VGND net130 sg13g2_tiehi
XFILLER_6_634 VPWR VGND sg13g2_fill_1
XFILLER_5_100 VPWR VGND sg13g2_fill_2
X_6553__169 VPWR VGND net169 sg13g2_tiehi
XFILLER_2_851 VPWR VGND sg13g2_decap_8
XFILLER_38_8 VPWR VGND sg13g2_fill_1
XFILLER_1_372 VPWR VGND sg13g2_fill_1
X_6685__570 VPWR VGND net754 sg13g2_tiehi
X_6761__480 VPWR VGND net664 sg13g2_tiehi
X_4870_ _1714_ _1709_ _1712_ VPWR VGND sg13g2_nand2b_1
XFILLER_32_210 VPWR VGND sg13g2_fill_1
X_3821_ _0772_ _0808_ _0859_ _0861_ VPWR VGND sg13g2_nor3_1
X_6460__274 VPWR VGND net274 sg13g2_tiehi
X_6540_ net182 VGND VPWR net1207 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[3\]
+ clknet_leaf_36_clk sg13g2_dfrbpq_1
X_6692__563 VPWR VGND net747 sg13g2_tiehi
X_3752_ _0800_ _0804_ _0805_ VPWR VGND sg13g2_and2_1
Xclkbuf_leaf_12_clk clknet_4_6_0_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
XFILLER_9_472 VPWR VGND sg13g2_fill_1
X_6471_ net253 VGND VPWR _0080_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[10\]
+ clknet_leaf_1_clk sg13g2_dfrbpq_1
X_3683_ _0720_ _0719_ _0736_ VPWR VGND sg13g2_xor2_1
X_5422_ _2162_ _2163_ _0315_ VPWR VGND sg13g2_nor2b_1
X_5353_ _2105_ _0557_ _2104_ VPWR VGND sg13g2_xnor2_1
X_4304_ _1241_ VPWR _1244_ VGND _0586_ net381 sg13g2_o21ai_1
X_5284_ _0293_ net496 _2046_ _2047_ VPWR VGND sg13g2_and3_1
X_4235_ _1185_ net1309 net383 VPWR VGND sg13g2_xnor2_1
X_4166_ _1126_ net1355 _1124_ VPWR VGND sg13g2_xnor2_1
X_4097_ _0080_ net441 _1071_ _1072_ VPWR VGND sg13g2_and3_1
X_6877__331 VPWR VGND net331 sg13g2_tiehi
X_6807_ net618 VGND VPWR _0416_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[2\]
+ clknet_leaf_62_clk sg13g2_dfrbpq_2
XFILLER_12_928 VPWR VGND sg13g2_decap_8
X_4999_ net426 _1820_ _1821_ _0234_ VPWR VGND sg13g2_nor3_1
X_6738_ net687 VGND VPWR _0347_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[9\]
+ clknet_leaf_56_clk sg13g2_dfrbpq_2
XFILLER_20_961 VPWR VGND sg13g2_decap_8
X_6669_ net53 VGND VPWR net1246 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[6\]\[3\]
+ clknet_leaf_51_clk sg13g2_dfrbpq_1
XFILLER_48_21 VPWR VGND sg13g2_decap_8
Xfanout440 _0546_ net440 VPWR VGND sg13g2_buf_8
Xfanout484 net485 net484 VPWR VGND sg13g2_buf_1
Xfanout451 net851 net451 VPWR VGND sg13g2_buf_8
Xfanout473 net851 net473 VPWR VGND sg13g2_buf_8
XFILLER_24_1023 VPWR VGND sg13g2_decap_4
Xfanout462 net466 net462 VPWR VGND sg13g2_buf_8
XFILLER_48_87 VPWR VGND sg13g2_decap_4
Xfanout495 net505 net495 VPWR VGND sg13g2_buf_1
XFILLER_11_961 VPWR VGND sg13g2_decap_8
XFILLER_7_932 VPWR VGND sg13g2_decap_8
XFILLER_31_1027 VPWR VGND sg13g2_fill_2
XFILLER_6_453 VPWR VGND sg13g2_fill_2
X_4020_ VGND VPWR _1012_ _1013_ _1016_ _1011_ sg13g2_a21oi_1
Xclkbuf_leaf_1_clk clknet_4_0_0_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
X_6529__193 VPWR VGND net193 sg13g2_tiehi
X_5971_ _2617_ VPWR _2627_ VGND _0581_ _2622_ sg13g2_o21ai_1
XFILLER_37_368 VPWR VGND sg13g2_fill_2
X_4922_ _1753_ VPWR _1758_ VGND _1754_ _1756_ sg13g2_o21ai_1
X_4853_ _1660_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[10\]
+ _1700_ VPWR VGND sg13g2_xor2_1
X_4784_ _1642_ net1365 _1640_ VPWR VGND sg13g2_xnor2_1
X_3804_ VGND VPWR net553 _0847_ _0012_ net883 sg13g2_a21oi_1
X_3735_ _0768_ _0787_ _0747_ _0788_ VPWR VGND sg13g2_nand3_1
X_6523_ net199 VGND VPWR net819 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].z_sign
+ clknet_leaf_42_clk sg13g2_dfrbpq_2
X_6454_ net285 VGND VPWR net886 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[7\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_2
X_6536__186 VPWR VGND net186 sg13g2_tiehi
X_5405_ net1054 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[4\] _2149_
+ VPWR VGND sg13g2_nor2b_1
X_3666_ _0719_ _0639_ _0699_ VPWR VGND sg13g2_xnor2_1
X_6385_ VGND VPWR net402 _2882_ _0467_ _2886_ sg13g2_a21oi_1
X_3597_ _0641_ net408 net404 net403 _0650_ VPWR VGND sg13g2_nor4_1
X_5336_ _2090_ net1255 _2088_ VPWR VGND sg13g2_xnor2_1
X_5267_ net489 net772 _0288_ VPWR VGND sg13g2_and2_1
X_4218_ net486 VPWR _1171_ VGND _1169_ _1170_ sg13g2_o21ai_1
X_6582__140 VPWR VGND net140 sg13g2_tiehi
X_5198_ VGND VPWR _0568_ _1969_ _1977_ net527 sg13g2_a21oi_1
X_4149_ VGND VPWR _1110_ _1111_ _0093_ _1112_ sg13g2_a21oi_1
X_6543__179 VPWR VGND net179 sg13g2_tiehi
XFILLER_34_34 VPWR VGND sg13g2_fill_1
Xclkload0 clknet_4_1_0_clk clkload0/X VPWR VGND sg13g2_buf_8
XFILLER_4_902 VPWR VGND sg13g2_decap_8
X_6751__490 VPWR VGND net674 sg13g2_tiehi
XFILLER_4_979 VPWR VGND sg13g2_decap_8
X_6897__548 VPWR VGND net732 sg13g2_tiehi
XFILLER_42_393 VPWR VGND sg13g2_fill_2
X_3520_ VPWR _0590_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[8\] VGND
+ sg13g2_inv_1
Xhold707 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[2\] VPWR VGND net1464
+ sg13g2_dlygate4sd3_1
Xhold718 _2485_ VPWR VGND net1475 sg13g2_dlygate4sd3_1
Xhold729 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[11\] VPWR VGND net1486
+ sg13g2_dlygate4sd3_1
X_6170_ VGND VPWR _2786_ _2790_ _2792_ net424 sg13g2_a21oi_1
XFILLER_3_990 VPWR VGND sg13g2_decap_8
X_5121_ _1912_ net1275 _1909_ VPWR VGND sg13g2_xnor2_1
X_5052_ _1850_ _1853_ _1864_ _1865_ VPWR VGND sg13g2_or3_1
X_4003_ _0997_ _1000_ _0994_ _1002_ VPWR VGND sg13g2_nand3_1
X_6661__61 VPWR VGND net61 sg13g2_tiehi
XFILLER_25_316 VPWR VGND sg13g2_fill_2
X_5954_ _2613_ _2608_ _2612_ VPWR VGND sg13g2_nand2_1
X_5885_ VGND VPWR _2551_ _2552_ _0388_ _2553_ sg13g2_a21oi_1
XFILLER_21_511 VPWR VGND sg13g2_fill_1
X_4905_ _1743_ _1731_ _1742_ VPWR VGND sg13g2_nand2_1
X_4836_ VGND VPWR net1137 net392 _1686_ _1683_ sg13g2_a21oi_1
XFILLER_14_1011 VPWR VGND sg13g2_decap_8
X_4767_ net488 VPWR _1628_ VGND _1626_ _1627_ sg13g2_o21ai_1
X_6506_ net216 VGND VPWR _0115_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[7\]
+ clknet_leaf_41_clk sg13g2_dfrbpq_2
X_3718_ VGND VPWR _0697_ _0765_ _0771_ _0764_ sg13g2_a21oi_1
X_4698_ _1566_ VPWR _1569_ VGND _1562_ _1567_ sg13g2_o21ai_1
X_6437_ net310 VGND VPWR _0046_ u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[3\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
X_3649_ _0700_ _0701_ _0702_ VPWR VGND sg13g2_nor2_1
X_6368_ net377 VPWR _2922_ VGND net1022 _2919_ sg13g2_o21ai_1
X_5319_ VGND VPWR _2075_ _2074_ _0554_ sg13g2_or2_1
XFILLER_1_938 VPWR VGND sg13g2_decap_8
X_6299_ _2872_ _2882_ _2893_ VPWR VGND sg13g2_nor2b_1
Xhold23 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[8\] VPWR VGND net780
+ sg13g2_dlygate4sd3_1
Xhold12 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[3\] VPWR VGND net769
+ sg13g2_dlygate4sd3_1
Xhold45 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[1\] VPWR VGND net802
+ sg13g2_dlygate4sd3_1
Xhold56 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[10\] VPWR VGND net813 sg13g2_dlygate4sd3_1
Xhold34 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[0\] VPWR VGND net791
+ sg13g2_dlygate4sd3_1
Xhold78 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[9\] VPWR VGND net835 sg13g2_dlygate4sd3_1
Xhold67 u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[5\] VPWR VGND net824 sg13g2_dlygate4sd3_1
Xhold89 u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[4\] VPWR VGND net846 sg13g2_dlygate4sd3_1
XFILLER_29_644 VPWR VGND sg13g2_fill_2
XFILLER_43_157 VPWR VGND sg13g2_fill_1
XFILLER_6_38 VPWR VGND sg13g2_fill_1
XFILLER_4_776 VPWR VGND sg13g2_decap_8
XFILLER_19_154 VPWR VGND sg13g2_fill_2
X_6526__196 VPWR VGND net196 sg13g2_tiehi
X_5670_ VGND VPWR net412 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[6\]
+ _2372_ _2365_ sg13g2_a21oi_1
X_4621_ VGND VPWR _1498_ _1503_ _1505_ net433 sg13g2_a21oi_1
X_4552_ _1449_ net760 _1448_ VPWR VGND sg13g2_nand2_1
X_6457__279 VPWR VGND net279 sg13g2_tiehi
X_6572__150 VPWR VGND net150 sg13g2_tiehi
Xhold515 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[2\] VPWR VGND net1272
+ sg13g2_dlygate4sd3_1
X_3503_ VPWR _0573_ net512 VGND sg13g2_inv_1
Xhold526 _0439_ VPWR VGND net1283 sg13g2_dlygate4sd3_1
X_4483_ VGND VPWR _1384_ _1390_ _1392_ net433 sg13g2_a21oi_1
Xhold504 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[1\] VPWR
+ VGND net1261 sg13g2_dlygate4sd3_1
Xhold537 _0189_ VPWR VGND net1294 sg13g2_dlygate4sd3_1
Xhold548 _0314_ VPWR VGND net1305 sg13g2_dlygate4sd3_1
Xhold559 _0287_ VPWR VGND net1316 sg13g2_dlygate4sd3_1
X_6222_ _2829_ _2827_ _2832_ _2834_ VPWR VGND sg13g2_a21o_1
X_6533__189 VPWR VGND net189 sg13g2_tiehi
XFILLER_44_1026 VPWR VGND sg13g2_fill_2
X_6153_ net453 VPWR _2777_ VGND _2771_ _2775_ sg13g2_o21ai_1
X_5104_ _1890_ _1896_ _1897_ VPWR VGND sg13g2_nor2_1
X_6084_ _0423_ net454 net1498 _2717_ VPWR VGND sg13g2_and3_1
X_5035_ _1850_ VPWR _1851_ VGND _0618_ net396 sg13g2_o21ai_1
XFILLER_39_986 VPWR VGND sg13g2_fill_2
X_5937_ _2598_ net1326 _2597_ VPWR VGND sg13g2_xnor2_1
X_6405__370 VPWR VGND net370 sg13g2_tiehi
X_5868_ VGND VPWR _2533_ _2537_ _2539_ _2536_ sg13g2_a21oi_1
X_5799_ _2477_ _2478_ _2479_ VPWR VGND sg13g2_nor2b_1
XFILLER_21_385 VPWR VGND sg13g2_fill_2
X_4819_ _1669_ _1671_ _1672_ VPWR VGND sg13g2_and2_1
XFILLER_1_735 VPWR VGND sg13g2_decap_8
XFILLER_44_455 VPWR VGND sg13g2_fill_1
XFILLER_12_330 VPWR VGND sg13g2_fill_2
XFILLER_13_853 VPWR VGND sg13g2_fill_1
XFILLER_12_341 VPWR VGND sg13g2_fill_2
XFILLER_39_216 VPWR VGND sg13g2_fill_1
X_6840_ net585 VGND VPWR net1073 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[9\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_35_444 VPWR VGND sg13g2_fill_2
XFILLER_36_989 VPWR VGND sg13g2_fill_1
X_6771_ net654 VGND VPWR net1349 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[4\]
+ clknet_leaf_60_clk sg13g2_dfrbpq_2
X_5722_ _2418_ net1549 _2416_ VPWR VGND sg13g2_xnor2_1
X_3983_ _0983_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[16\] _0984_
+ VPWR VGND sg13g2_nor2b_2
X_5653_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[3\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[4\]
+ _2357_ VPWR VGND sg13g2_nor2_1
X_4604_ VGND VPWR _0608_ net832 _0170_ _1490_ sg13g2_a21oi_1
X_5584_ net474 VPWR _2299_ VGND _2293_ _2298_ sg13g2_o21ai_1
XFILLER_11_1003 VPWR VGND sg13g2_decap_8
X_6394__388 VPWR VGND net572 sg13g2_tiehi
Xhold301 _1079_ VPWR VGND net1058 sg13g2_dlygate4sd3_1
X_4535_ _1436_ _1433_ _1434_ _1435_ VPWR VGND sg13g2_and3_1
Xhold312 _2651_ VPWR VGND net1069 sg13g2_dlygate4sd3_1
Xhold334 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[6\] VPWR VGND net1091
+ sg13g2_dlygate4sd3_1
Xhold323 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[4\] VPWR VGND net1080
+ sg13g2_dlygate4sd3_1
Xhold345 _0263_ VPWR VGND net1102 sg13g2_dlygate4sd3_1
Xhold367 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[8\] VPWR VGND net1124
+ sg13g2_dlygate4sd3_1
X_4466_ _1377_ net985 net996 VPWR VGND sg13g2_nand2_1
Xhold356 _0229_ VPWR VGND net1113 sg13g2_dlygate4sd3_1
Xhold378 _1476_ VPWR VGND net1135 sg13g2_dlygate4sd3_1
Xhold389 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[2\]\[1\] VPWR VGND net1146
+ sg13g2_dlygate4sd3_1
X_6205_ net508 net1005 _2820_ VPWR VGND sg13g2_xor2_1
X_4397_ VGND VPWR _1311_ _1317_ _1319_ net436 sg13g2_a21oi_1
X_6136_ _2757_ net1547 _2762_ VPWR VGND sg13g2_nor2_1
X_6067_ _2691_ _2695_ _2702_ _2703_ VPWR VGND sg13g2_nor3_1
X_5018_ _1836_ net1488 _1837_ VPWR VGND sg13g2_nor2b_1
XFILLER_14_639 VPWR VGND sg13g2_fill_1
XFILLER_13_149 VPWR VGND sg13g2_fill_1
XFILLER_21_160 VPWR VGND sg13g2_fill_1
XFILLER_18_912 VPWR VGND sg13g2_decap_8
X_6562__160 VPWR VGND net160 sg13g2_tiehi
XFILLER_45_764 VPWR VGND sg13g2_fill_2
XFILLER_18_989 VPWR VGND sg13g2_decap_8
X_6523__199 VPWR VGND net199 sg13g2_tiehi
X_4320_ _1255_ _1256_ _1248_ _1257_ VPWR VGND sg13g2_nand3_1
X_4251_ _1196_ net1277 _1198_ VPWR VGND sg13g2_xor2_1
X_4182_ _1139_ net1499 _1140_ VPWR VGND sg13g2_nor2b_1
XFILLER_27_219 VPWR VGND sg13g2_fill_1
X_6823_ net602 VGND VPWR net1407 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[3\]
+ clknet_leaf_60_clk sg13g2_dfrbpq_2
X_6754_ net671 VGND VPWR net905 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[10\]
+ clknet_leaf_57_clk sg13g2_dfrbpq_2
X_3966_ _0967_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[7\] _0945_
+ VPWR VGND sg13g2_xnor2_1
X_5705_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[5\] _2402_
+ _2403_ VPWR VGND sg13g2_and2_1
X_6685_ net754 VGND VPWR net1145 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[6\]
+ clknet_leaf_44_clk sg13g2_dfrbpq_1
X_3897_ VGND VPWR u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[5\] _0915_ _0917_ net941
+ sg13g2_a21oi_1
X_5636_ _2344_ net1194 _2336_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_808 VPWR VGND sg13g2_decap_8
X_5567_ VGND VPWR _2277_ _2282_ _0340_ _2283_ sg13g2_a21oi_1
X_4518_ net1537 net384 _1422_ VPWR VGND sg13g2_nor2_1
Xhold131 _0893_ VPWR VGND net888 sg13g2_dlygate4sd3_1
Xhold153 _0853_ VPWR VGND net910 sg13g2_dlygate4sd3_1
Xhold142 _2900_ VPWR VGND net899 sg13g2_dlygate4sd3_1
Xhold120 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[1\] VPWR VGND net877
+ sg13g2_dlygate4sd3_1
X_5498_ net482 VPWR _2228_ VGND net852 _2227_ sg13g2_o21ai_1
Xhold164 _0033_ VPWR VGND net921 sg13g2_dlygate4sd3_1
Xhold186 _0037_ VPWR VGND net943 sg13g2_dlygate4sd3_1
Xhold175 _2902_ VPWR VGND net932 sg13g2_dlygate4sd3_1
X_4449_ _1361_ net1370 _1363_ VPWR VGND sg13g2_nor2b_1
Xhold197 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[3\] VPWR VGND
+ net954 sg13g2_dlygate4sd3_1
X_6847__394 VPWR VGND net578 sg13g2_tiehi
X_6119_ VGND VPWR _2747_ _2745_ net1552 sg13g2_or2_1
XFILLER_2_1012 VPWR VGND sg13g2_decap_8
XFILLER_27_764 VPWR VGND sg13g2_fill_2
XFILLER_15_948 VPWR VGND sg13g2_decap_8
XFILLER_23_992 VPWR VGND sg13g2_decap_8
XFILLER_10_653 VPWR VGND sg13g2_fill_1
XFILLER_5_134 VPWR VGND sg13g2_fill_2
XFILLER_2_830 VPWR VGND sg13g2_decap_8
X_6677__45 VPWR VGND net45 sg13g2_tiehi
XFILLER_17_252 VPWR VGND sg13g2_fill_2
XFILLER_32_200 VPWR VGND sg13g2_fill_2
X_3820_ _0858_ VPWR _0860_ VGND _0809_ _0859_ sg13g2_o21ai_1
X_3751_ _0801_ net403 _0804_ VPWR VGND sg13g2_xor2_1
X_6470_ net255 VGND VPWR _0079_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[9\]
+ clknet_leaf_1_clk sg13g2_dfrbpq_2
X_3682_ _0730_ _0731_ _0725_ _0735_ VPWR VGND sg13g2_nand3_1
X_5421_ VGND VPWR _2156_ _2161_ _2163_ net429 sg13g2_a21oi_1
X_5352_ net521 _2094_ _2104_ VPWR VGND sg13g2_nor2_1
X_4303_ VPWR _1243_ _1242_ VGND sg13g2_inv_1
X_5283_ _2042_ _2040_ _2045_ _2047_ VPWR VGND sg13g2_a21o_1
X_4234_ _1181_ _1183_ _1184_ VPWR VGND sg13g2_nor2_1
X_4165_ _1124_ net1355 _1125_ VPWR VGND sg13g2_nor2b_1
X_4096_ net865 _1069_ net859 _1072_ VPWR VGND sg13g2_nand3_1
X_6806_ net619 VGND VPWR net1077 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[1\]
+ clknet_leaf_62_clk sg13g2_dfrbpq_1
XFILLER_12_907 VPWR VGND sg13g2_decap_8
XFILLER_11_428 VPWR VGND sg13g2_fill_2
XFILLER_23_277 VPWR VGND sg13g2_fill_1
X_4998_ VGND VPWR _1815_ _1819_ _1821_ _1818_ sg13g2_a21oi_1
X_6737_ net688 VGND VPWR net1336 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[8\]
+ clknet_leaf_55_clk sg13g2_dfrbpq_1
XFILLER_20_940 VPWR VGND sg13g2_decap_8
X_3949_ _0950_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[13\] _0949_
+ VPWR VGND sg13g2_xnor2_1
X_6668_ net54 VGND VPWR _0277_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[6\]\[2\]
+ clknet_leaf_51_clk sg13g2_dfrbpq_1
X_5619_ VGND VPWR _0597_ _2321_ _2329_ net516 sg13g2_a21oi_1
X_6599_ net123 VGND VPWR _0208_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].y_shr\[0\]
+ clknet_leaf_27_clk sg13g2_dfrbpq_2
X_6552__170 VPWR VGND net170 sg13g2_tiehi
Xfanout441 net443 net441 VPWR VGND sg13g2_buf_8
Xfanout430 net434 net430 VPWR VGND sg13g2_buf_2
X_6674__48 VPWR VGND net48 sg13g2_tiehi
XFILLER_24_1002 VPWR VGND sg13g2_decap_8
Xfanout463 net465 net463 VPWR VGND sg13g2_buf_2
Xfanout452 net456 net452 VPWR VGND sg13g2_buf_8
Xfanout474 net476 net474 VPWR VGND sg13g2_buf_8
XFILLER_48_77 VPWR VGND sg13g2_decap_4
Xfanout485 net490 net485 VPWR VGND sg13g2_buf_8
Xfanout496 net500 net496 VPWR VGND sg13g2_buf_8
XFILLER_27_550 VPWR VGND sg13g2_fill_1
XFILLER_15_756 VPWR VGND sg13g2_fill_2
XFILLER_42_597 VPWR VGND sg13g2_fill_1
XFILLER_11_940 VPWR VGND sg13g2_decap_8
XFILLER_7_911 VPWR VGND sg13g2_decap_8
XFILLER_7_988 VPWR VGND sg13g2_decap_8
X_5970_ net425 _2625_ _2626_ _0400_ VPWR VGND sg13g2_nor3_1
X_4921_ _1753_ _1754_ _1756_ _1757_ VPWR VGND sg13g2_nor3_1
X_4852_ _1697_ net1202 _1691_ _1699_ VPWR VGND sg13g2_nand3_1
X_3803_ net553 net882 _0848_ VPWR VGND sg13g2_nor2_1
X_4783_ _1641_ net1365 _1640_ VPWR VGND sg13g2_nand2_1
X_3734_ _0787_ _0772_ _0786_ VPWR VGND sg13g2_xnor2_1
X_6522_ net200 VGND VPWR _0131_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[10\]
+ clknet_leaf_42_clk sg13g2_dfrbpq_1
X_3665_ _0718_ _0640_ net406 VPWR VGND sg13g2_nand2_1
X_6453_ net287 VGND VPWR net953 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[6\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_2
X_5404_ VGND VPWR _2146_ _2147_ _0312_ _2148_ sg13g2_a21oi_1
X_6384_ _2879_ _2868_ _0464_ VPWR VGND sg13g2_nor2b_1
X_3596_ _0638_ _0640_ net407 net406 _0649_ VPWR VGND sg13g2_nor4_1
X_5335_ _2089_ net1255 _2088_ VPWR VGND sg13g2_nand2_1
X_5266_ VGND VPWR net1315 _2034_ _0287_ _2035_ sg13g2_a21oi_1
X_4217_ VGND VPWR net1183 net382 _1170_ _1167_ sg13g2_a21oi_1
X_6844__397 VPWR VGND net581 sg13g2_tiehi
X_5197_ VGND VPWR _1968_ _1973_ _1976_ _1972_ sg13g2_a21oi_1
X_4148_ net501 VPWR _1112_ VGND _1110_ _1111_ sg13g2_o21ai_1
X_4079_ _1059_ net846 _1061_ VPWR VGND sg13g2_xor2_1
Xclkload1 clknet_4_2_0_clk clkload1/X VPWR VGND sg13g2_buf_8
XFILLER_4_958 VPWR VGND sg13g2_decap_8
X_6415__350 VPWR VGND net350 sg13g2_tiehi
XFILLER_46_199 VPWR VGND sg13g2_fill_2
XFILLER_43_884 VPWR VGND sg13g2_fill_2
XFILLER_30_501 VPWR VGND sg13g2_decap_8
Xhold708 _1786_ VPWR VGND net1465 sg13g2_dlygate4sd3_1
XFILLER_7_785 VPWR VGND sg13g2_fill_2
Xhold719 _0379_ VPWR VGND net1476 sg13g2_dlygate4sd3_1
X_5120_ VPWR _1911_ _1910_ VGND sg13g2_inv_1
X_5051_ _1858_ VPWR _1864_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[7\]
+ net395 sg13g2_o21ai_1
X_4002_ VGND VPWR _0994_ _0997_ _1001_ _1000_ sg13g2_a21oi_1
XFILLER_26_807 VPWR VGND sg13g2_fill_2
X_6542__180 VPWR VGND net180 sg13g2_tiehi
X_5953_ _2610_ net1457 _2612_ VPWR VGND sg13g2_xor2_1
X_4904_ net389 VPWR _1742_ VGND net1432 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[7\]
+ sg13g2_o21ai_1
X_5884_ net459 VPWR _2553_ VGND _2551_ _2552_ sg13g2_o21ai_1
X_4835_ VPWR _1685_ _1684_ VGND sg13g2_inv_1
X_4766_ net401 net1399 _1627_ VPWR VGND sg13g2_xor2_1
X_6505_ net217 VGND VPWR _0114_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[6\]
+ clknet_leaf_36_clk sg13g2_dfrbpq_1
X_3717_ _0698_ _0766_ _0770_ VPWR VGND sg13g2_nor2_1
X_4697_ VGND VPWR _1562_ _1567_ _0185_ _1568_ sg13g2_a21oi_1
X_6436_ net311 VGND VPWR _0045_ u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[2\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
X_3648_ _0701_ _0637_ _0653_ VPWR VGND sg13g2_xnor2_1
X_3579_ _0635_ net859 u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[11\] VPWR VGND
+ sg13g2_nand2b_1
XFILLER_1_917 VPWR VGND sg13g2_decap_8
X_6367_ net1022 _2919_ _2921_ VPWR VGND sg13g2_and2_1
X_5318_ _2074_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[1\]
+ _2073_ VPWR VGND sg13g2_xnor2_1
Xhold13 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[0\] VPWR VGND net770
+ sg13g2_dlygate4sd3_1
X_6298_ _0471_ net444 _2891_ _2892_ VPWR VGND sg13g2_and3_1
Xhold24 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[6\] VPWR VGND net781
+ sg13g2_dlygate4sd3_1
Xhold35 u_angle_cordic_12b_pmod.u_vga_top.clk_div_cnt\[0\] VPWR VGND net792 sg13g2_dlygate4sd3_1
X_5249_ VGND VPWR _2019_ _2020_ _0284_ _2021_ sg13g2_a21oi_1
Xhold46 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[11\] VPWR VGND
+ net803 sg13g2_dlygate4sd3_1
Xhold68 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[11\] VPWR VGND net825
+ sg13g2_dlygate4sd3_1
Xhold57 _0006_ VPWR VGND net814 sg13g2_dlygate4sd3_1
Xhold79 _0005_ VPWR VGND net836 sg13g2_dlygate4sd3_1
XFILLER_45_34 VPWR VGND sg13g2_fill_2
XFILLER_24_383 VPWR VGND sg13g2_fill_1
XFILLER_4_755 VPWR VGND sg13g2_decap_8
XFILLER_0_983 VPWR VGND sg13g2_decap_8
XFILLER_37_1001 VPWR VGND sg13g2_fill_2
X_4620_ _1498_ _1503_ _1504_ VPWR VGND sg13g2_nor2_1
X_4551_ net1006 net539 _1448_ VPWR VGND sg13g2_xor2_1
Xhold516 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[10\] VPWR VGND net1273
+ sg13g2_dlygate4sd3_1
X_3502_ VPWR _0572_ net1259 VGND sg13g2_inv_1
X_4482_ _1384_ net1224 _1391_ VPWR VGND sg13g2_nor2_1
Xhold505 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[12\] VPWR VGND net1262
+ sg13g2_dlygate4sd3_1
Xhold527 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[3\] VPWR VGND net1284
+ sg13g2_dlygate4sd3_1
Xhold549 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[6\] VPWR VGND net1306
+ sg13g2_dlygate4sd3_1
Xhold538 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[4\] VPWR VGND net1295
+ sg13g2_dlygate4sd3_1
X_6221_ _2829_ _2832_ _2827_ _2833_ VPWR VGND sg13g2_nand3_1
X_6152_ VPWR _2776_ _2775_ VGND sg13g2_inv_1
X_5103_ _1894_ net1393 _1896_ VPWR VGND sg13g2_xor2_1
XFILLER_32_0 VPWR VGND sg13g2_fill_2
X_6083_ _2711_ _2708_ _2715_ _2717_ VPWR VGND sg13g2_a21o_1
X_5034_ _0240_ net470 _1849_ _1850_ VPWR VGND sg13g2_and3_1
XFILLER_25_103 VPWR VGND sg13g2_fill_2
X_5936_ _2590_ VPWR _2597_ VGND net514 _0580_ sg13g2_o21ai_1
X_6737__504 VPWR VGND net688 sg13g2_tiehi
X_5867_ VGND VPWR _2533_ net1327 _0385_ _2538_ sg13g2_a21oi_1
X_5798_ _2478_ _0574_ _2476_ VPWR VGND sg13g2_nand2_1
XFILLER_31_14 VPWR VGND sg13g2_fill_1
X_4818_ VPWR _1671_ _1670_ VGND sg13g2_inv_1
X_4749_ net401 net1504 _1613_ VPWR VGND sg13g2_xor2_1
X_6419_ net342 VGND VPWR net843 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[8\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_2
XFILLER_1_714 VPWR VGND sg13g2_decap_8
XFILLER_49_707 VPWR VGND sg13g2_fill_2
XFILLER_0_213 VPWR VGND sg13g2_fill_1
XFILLER_5_1010 VPWR VGND sg13g2_decap_8
XFILLER_9_869 VPWR VGND sg13g2_decap_8
X_6532__190 VPWR VGND net190 sg13g2_tiehi
XFILLER_0_780 VPWR VGND sg13g2_decap_8
XFILLER_48_740 VPWR VGND sg13g2_fill_1
X_6770_ net655 VGND VPWR net1476 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[3\]
+ clknet_leaf_61_clk sg13g2_dfrbpq_2
X_3982_ _0983_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[11\] _0948_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_44_990 VPWR VGND sg13g2_fill_2
X_5721_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[7\] _2416_
+ _2417_ VPWR VGND sg13g2_and2_1
X_5652_ _2353_ VPWR _2356_ VGND _2349_ _2354_ sg13g2_o21ai_1
XFILLER_30_150 VPWR VGND sg13g2_fill_1
X_5583_ _2298_ net1415 _2296_ VPWR VGND sg13g2_xnor2_1
X_4603_ VGND VPWR _1488_ _1489_ _0169_ _1490_ sg13g2_a21oi_1
Xhold302 _0086_ VPWR VGND net1059 sg13g2_dlygate4sd3_1
X_4534_ _1435_ net1169 net385 VPWR VGND sg13g2_xnor2_1
Xhold313 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[0\].y_shr\[11\] VPWR
+ VGND net1070 sg13g2_dlygate4sd3_1
Xhold335 _0205_ VPWR VGND net1092 sg13g2_dlygate4sd3_1
Xhold324 _0125_ VPWR VGND net1081 sg13g2_dlygate4sd3_1
X_6470__255 VPWR VGND net255 sg13g2_tiehi
Xhold346 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[6\]\[0\] VPWR VGND net1103
+ sg13g2_dlygate4sd3_1
Xhold357 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[6\] VPWR VGND net1114
+ sg13g2_dlygate4sd3_1
Xhold368 _2265_ VPWR VGND net1125 sg13g2_dlygate4sd3_1
X_4465_ VGND VPWR _1374_ _1375_ _0145_ _1376_ sg13g2_a21oi_1
X_4396_ _1311_ _1317_ _1318_ VPWR VGND sg13g2_nor2_1
X_6204_ _2819_ net1005 net508 VPWR VGND sg13g2_nand2_1
Xhold379 _0166_ VPWR VGND net1136 sg13g2_dlygate4sd3_1
X_6135_ _2761_ _0620_ _2759_ VPWR VGND sg13g2_xnor2_1
X_6066_ VPWR _2702_ _2701_ VGND sg13g2_inv_1
X_5017_ _1834_ _1835_ _1836_ VPWR VGND sg13g2_nor2b_1
XFILLER_26_434 VPWR VGND sg13g2_fill_2
X_5919_ _2578_ VPWR _2582_ VGND _2574_ _2579_ sg13g2_o21ai_1
X_6899_ net734 VGND VPWR _0527_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[6\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_6_839 VPWR VGND sg13g2_decap_8
XFILLER_18_968 VPWR VGND sg13g2_decap_8
XFILLER_29_294 VPWR VGND sg13g2_fill_2
XFILLER_33_949 VPWR VGND sg13g2_fill_1
XFILLER_8_165 VPWR VGND sg13g2_fill_1
XFILLER_4_382 VPWR VGND sg13g2_fill_2
X_4250_ net1277 _1196_ _1197_ VPWR VGND sg13g2_and2_1
X_4181_ _1137_ _1138_ _1139_ VPWR VGND sg13g2_nor2b_1
X_6727__514 VPWR VGND net698 sg13g2_tiehi
X_6822_ net603 VGND VPWR _0431_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[2\]
+ clknet_leaf_63_clk sg13g2_dfrbpq_2
XFILLER_17_990 VPWR VGND sg13g2_decap_8
X_6753_ net672 VGND VPWR net1119 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[7\]
+ clknet_leaf_57_clk sg13g2_dfrbpq_1
X_3965_ _0966_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[6\] _0965_
+ VPWR VGND sg13g2_xnor2_1
X_6734__507 VPWR VGND net691 sg13g2_tiehi
X_3896_ net420 _0916_ _0036_ VPWR VGND sg13g2_nor2_1
X_5704_ _2402_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[11\] _2401_
+ VPWR VGND sg13g2_xnor2_1
X_6684_ net755 VGND VPWR _0293_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[5\]
+ clknet_leaf_41_clk sg13g2_dfrbpq_1
X_5635_ _2336_ net1194 _2343_ VPWR VGND sg13g2_nor2b_1
XFILLER_31_481 VPWR VGND sg13g2_fill_1
X_5566_ net474 VPWR _2283_ VGND _2277_ _2282_ sg13g2_o21ai_1
Xhold110 _0857_ VPWR VGND net867 sg13g2_dlygate4sd3_1
X_4517_ VGND VPWR _1415_ _1418_ _1421_ _1417_ sg13g2_a21oi_1
Xhold121 u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[11\] VPWR VGND net878 sg13g2_dlygate4sd3_1
Xhold132 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[8\] VPWR VGND net889 sg13g2_dlygate4sd3_1
Xhold143 _0503_ VPWR VGND net900 sg13g2_dlygate4sd3_1
X_5497_ _2227_ net524 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[1\]
+ VPWR VGND sg13g2_xnor2_1
Xhold165 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[0\] VPWR VGND net922
+ sg13g2_dlygate4sd3_1
Xhold176 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[0\] VPWR VGND net933
+ sg13g2_dlygate4sd3_1
Xhold154 _0015_ VPWR VGND net911 sg13g2_dlygate4sd3_1
X_4448_ net386 VPWR _1362_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[1\]
+ net1369 sg13g2_o21ai_1
Xhold198 _0059_ VPWR VGND net955 sg13g2_dlygate4sd3_1
Xhold187 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[4\] VPWR VGND net944 sg13g2_dlygate4sd3_1
X_4379_ VGND VPWR net410 net818 _0132_ _1303_ sg13g2_a21oi_1
X_6118_ net1552 _2745_ _2746_ VPWR VGND sg13g2_and2_1
XFILLER_46_529 VPWR VGND sg13g2_fill_1
X_6049_ _2687_ net1209 _2685_ VPWR VGND sg13g2_xnor2_1
XFILLER_39_592 VPWR VGND sg13g2_fill_2
XFILLER_15_927 VPWR VGND sg13g2_decap_8
XFILLER_14_437 VPWR VGND sg13g2_fill_2
XFILLER_14_448 VPWR VGND sg13g2_fill_2
XFILLER_23_971 VPWR VGND sg13g2_decap_8
XFILLER_41_267 VPWR VGND sg13g2_fill_2
XFILLER_2_886 VPWR VGND sg13g2_decap_8
X_6425__330 VPWR VGND net330 sg13g2_tiehi
X_3750_ VPWR _0803_ _0802_ VGND sg13g2_inv_1
X_3681_ _0734_ _0731_ _0732_ VPWR VGND sg13g2_xnor2_1
X_5420_ _2156_ _2161_ _2162_ VPWR VGND sg13g2_nor2_1
X_5351_ VGND VPWR _2092_ _2099_ _2103_ _2098_ sg13g2_a21oi_1
X_4302_ net381 net1512 _1242_ VPWR VGND sg13g2_xor2_1
X_5282_ _2042_ _2045_ _2040_ _2046_ VPWR VGND sg13g2_nand3_1
X_4233_ _1183_ _1174_ _1182_ VPWR VGND sg13g2_nand2_1
X_4164_ _1124_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[8\] _1123_
+ VPWR VGND sg13g2_xnor2_1
X_4095_ _1069_ net865 net859 _1071_ VPWR VGND sg13g2_a21o_1
X_6805_ net620 VGND VPWR net1048 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[0\]
+ clknet_leaf_62_clk sg13g2_dfrbpq_1
X_6736_ net689 VGND VPWR net1403 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[7\]
+ clknet_leaf_55_clk sg13g2_dfrbpq_2
X_4997_ _1820_ _1815_ _1818_ _1819_ VPWR VGND sg13g2_and3_1
X_3948_ _0946_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[8\] _0949_
+ VPWR VGND sg13g2_xor2_1
X_6667_ net55 VGND VPWR net1064 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[6\]\[1\]
+ clknet_leaf_51_clk sg13g2_dfrbpq_1
X_3879_ _0904_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[1\] net1577 VPWR VGND sg13g2_nand2_1
X_5618_ _2325_ _2320_ _2324_ _2328_ VPWR VGND sg13g2_a21o_1
XFILLER_20_996 VPWR VGND sg13g2_decap_8
X_6598_ net124 VGND VPWR _0207_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[9\]
+ clknet_leaf_26_clk sg13g2_dfrbpq_2
X_5549_ net933 net1230 _2268_ VPWR VGND sg13g2_and2_1
Xfanout420 net423 net420 VPWR VGND sg13g2_buf_8
Xfanout431 net434 net431 VPWR VGND sg13g2_buf_8
Xfanout464 net465 net464 VPWR VGND sg13g2_buf_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
Xfanout453 net456 net453 VPWR VGND sg13g2_buf_1
Xfanout475 net476 net475 VPWR VGND sg13g2_buf_1
Xfanout442 net443 net442 VPWR VGND sg13g2_buf_1
Xfanout486 net487 net486 VPWR VGND sg13g2_buf_8
Xfanout497 net500 net497 VPWR VGND sg13g2_buf_1
XFILLER_46_348 VPWR VGND sg13g2_fill_1
XFILLER_30_716 VPWR VGND sg13g2_fill_2
X_6717__524 VPWR VGND net708 sg13g2_tiehi
XFILLER_7_967 VPWR VGND sg13g2_decap_8
XFILLER_11_996 VPWR VGND sg13g2_decap_8
XFILLER_2_683 VPWR VGND sg13g2_decap_8
X_6724__517 VPWR VGND net701 sg13g2_tiehi
X_4920_ VPWR _1756_ _1755_ VGND sg13g2_inv_1
X_4851_ net392 VPWR _1698_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[1\]
+ net1201 sg13g2_o21ai_1
X_3802_ _0847_ _0652_ _0746_ VPWR VGND sg13g2_xnor2_1
X_4782_ _1640_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[10\] _1639_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_14_790 VPWR VGND sg13g2_fill_1
X_3733_ _0786_ _0773_ _0784_ VPWR VGND sg13g2_xnor2_1
X_6521_ net201 VGND VPWR _0130_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[9\]
+ clknet_leaf_42_clk sg13g2_dfrbpq_1
X_3664_ _0717_ _0707_ _0708_ VPWR VGND sg13g2_xnor2_1
X_6452_ net289 VGND VPWR _0061_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[5\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_2
X_5403_ net479 VPWR _2148_ VGND _2146_ _2147_ sg13g2_o21ai_1
X_6383_ net422 _2873_ _2880_ _0463_ VPWR VGND sg13g2_nor3_1
X_3595_ VGND VPWR _0648_ _0639_ _0637_ sg13g2_or2_1
X_5334_ _2087_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[3\]
+ _2088_ VPWR VGND sg13g2_xor2_1
X_5265_ net492 VPWR _2035_ VGND _2033_ _2034_ sg13g2_o21ai_1
X_5196_ _1974_ _1975_ _0277_ VPWR VGND sg13g2_nor2b_1
X_4216_ _1169_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[3\]
+ net382 VPWR VGND sg13g2_xnor2_1
XFILLER_29_827 VPWR VGND sg13g2_fill_2
X_4147_ _1111_ net533 net1036 VPWR VGND sg13g2_xnor2_1
X_4078_ net445 _1060_ _0073_ VPWR VGND sg13g2_and2_1
Xclkload2 clknet_4_3_0_clk clkload2/X VPWR VGND sg13g2_buf_8
X_6719_ net706 VGND VPWR net1075 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[2\]
+ clknet_leaf_31_clk sg13g2_dfrbpq_2
XFILLER_4_937 VPWR VGND sg13g2_decap_8
XFILLER_19_348 VPWR VGND sg13g2_fill_2
XFILLER_46_134 VPWR VGND sg13g2_fill_2
X_6670__52 VPWR VGND net52 sg13g2_tiehi
Xhold709 _0227_ VPWR VGND net1466 sg13g2_dlygate4sd3_1
XFILLER_7_775 VPWR VGND sg13g2_fill_2
XFILLER_7_753 VPWR VGND sg13g2_decap_8
X_5050_ VGND VPWR _1861_ _1862_ _0243_ _1863_ sg13g2_a21oi_1
X_4001_ _1000_ net980 net550 VPWR VGND sg13g2_xnor2_1
XFILLER_37_134 VPWR VGND sg13g2_fill_1
X_5952_ _2611_ net1457 _2610_ VPWR VGND sg13g2_nand2_1
X_4903_ _1721_ _1723_ _1728_ _1740_ _1741_ VPWR VGND sg13g2_nor4_1
X_5883_ _2552_ net1217 _2547_ VPWR VGND sg13g2_xnor2_1
X_4834_ _1684_ net1044 _1660_ VPWR VGND sg13g2_xnor2_1
X_4765_ _1625_ VPWR _1626_ VGND _1616_ _1624_ sg13g2_o21ai_1
X_3716_ _0769_ _0747_ _0768_ VPWR VGND sg13g2_nand2_1
X_6504_ net218 VGND VPWR net1405 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[5\]
+ clknet_leaf_36_clk sg13g2_dfrbpq_1
X_4696_ net482 VPWR _1568_ VGND _1562_ _1567_ sg13g2_o21ai_1
X_6850__391 VPWR VGND net575 sg13g2_tiehi
X_3647_ _0700_ _0639_ _0699_ VPWR VGND sg13g2_nand2_1
X_6435_ net312 VGND VPWR _0044_ u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[1\]
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
X_3578_ _0633_ _0634_ _0000_ VPWR VGND sg13g2_nor2_1
X_6366_ net375 _2919_ net959 _0514_ VPWR VGND sg13g2_nor3_1
X_5317_ net521 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[0\]
+ _2073_ VPWR VGND sg13g2_nor2b_1
X_6297_ _2889_ _2870_ _2883_ _2892_ VPWR VGND sg13g2_a21o_1
Xhold14 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[6\] VPWR VGND net771
+ sg13g2_dlygate4sd3_1
Xhold25 _0049_ VPWR VGND net782 sg13g2_dlygate4sd3_1
X_5248_ net480 VPWR _2021_ VGND _2019_ _2020_ sg13g2_o21ai_1
XFILLER_29_36 VPWR VGND sg13g2_fill_2
Xhold47 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[2\] VPWR VGND net804
+ sg13g2_dlygate4sd3_1
Xhold36 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[4\] VPWR VGND net793
+ sg13g2_dlygate4sd3_1
Xhold58 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[10\] VPWR VGND net815
+ sg13g2_dlygate4sd3_1
X_5179_ net912 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[5\] _1961_
+ VPWR VGND sg13g2_nor2b_1
X_6707__534 VPWR VGND net718 sg13g2_tiehi
XFILLER_21_1017 VPWR VGND sg13g2_decap_8
Xhold69 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[10\] VPWR VGND net826
+ sg13g2_dlygate4sd3_1
XFILLER_29_646 VPWR VGND sg13g2_fill_1
XFILLER_21_1028 VPWR VGND sg13g2_fill_1
X_6714__527 VPWR VGND net711 sg13g2_tiehi
XFILLER_4_734 VPWR VGND sg13g2_decap_8
XFILLER_0_962 VPWR VGND sg13g2_decap_8
XFILLER_19_145 VPWR VGND sg13g2_fill_1
XFILLER_19_156 VPWR VGND sg13g2_fill_1
XFILLER_28_690 VPWR VGND sg13g2_fill_1
X_4550_ _1447_ net539 net1006 VPWR VGND sg13g2_nand2_1
Xhold517 _0195_ VPWR VGND net1274 sg13g2_dlygate4sd3_1
X_3501_ _0571_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[10\] VPWR VGND
+ sg13g2_inv_2
X_4481_ _1388_ net1223 _1390_ VPWR VGND sg13g2_xor2_1
Xhold506 _0158_ VPWR VGND net1263 sg13g2_dlygate4sd3_1
Xhold539 _2680_ VPWR VGND net1296 sg13g2_dlygate4sd3_1
Xhold528 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[10\] VPWR
+ VGND net1285 sg13g2_dlygate4sd3_1
X_6220_ _2832_ net509 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[5\]
+ VPWR VGND sg13g2_xnor2_1
X_6151_ _2775_ net1420 _2773_ VPWR VGND sg13g2_xnor2_1
XFILLER_44_1028 VPWR VGND sg13g2_fill_1
X_5102_ net1393 _1894_ _1895_ VPWR VGND sg13g2_and2_1
X_6082_ _2711_ _2715_ _2708_ _2716_ VPWR VGND sg13g2_nand3_1
XFILLER_25_0 VPWR VGND sg13g2_fill_2
X_5033_ _1847_ _1844_ _1848_ _1850_ VPWR VGND sg13g2_a21o_2
X_5935_ _2593_ _2589_ _2592_ _2596_ VPWR VGND sg13g2_a21o_1
X_5866_ net459 VPWR _2538_ VGND _2533_ _2537_ sg13g2_o21ai_1
Xclkbuf_leaf_60_clk clknet_4_2_0_clk clknet_leaf_60_clk VPWR VGND sg13g2_buf_8
X_4817_ _1670_ net1091 net391 VPWR VGND sg13g2_xnor2_1
X_5797_ _0574_ _2476_ _2477_ VPWR VGND sg13g2_nor2_1
X_4748_ net400 net1526 _1610_ _1612_ VPWR VGND sg13g2_a21o_1
X_4679_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[3\] _1523_
+ _1554_ VPWR VGND sg13g2_and2_1
X_6418_ net344 VGND VPWR net1021 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[7\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_2
X_6349_ net374 _2908_ net1108 _0508_ VPWR VGND sg13g2_nor3_1
XFILLER_16_148 VPWR VGND sg13g2_fill_2
XFILLER_13_833 VPWR VGND sg13g2_fill_1
XFILLER_12_343 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_51_clk clknet_4_10_0_clk clknet_leaf_51_clk VPWR VGND sg13g2_buf_8
XFILLER_9_848 VPWR VGND sg13g2_decap_8
XFILLER_13_888 VPWR VGND sg13g2_decap_8
X_6456__281 VPWR VGND net281 sg13g2_tiehi
X_6864__357 VPWR VGND net357 sg13g2_tiehi
XFILLER_47_284 VPWR VGND sg13g2_fill_2
X_3981_ _0982_ _0979_ _0981_ VPWR VGND sg13g2_nand2_1
X_5720_ VGND VPWR _2410_ _2416_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[12\]
+ net520 sg13g2_a21oi_2
Xclkbuf_leaf_42_clk clknet_4_14_0_clk clknet_leaf_42_clk VPWR VGND sg13g2_buf_8
X_5651_ VGND VPWR _2349_ _2354_ _0352_ _2355_ sg13g2_a21oi_1
XFILLER_31_674 VPWR VGND sg13g2_fill_2
X_4602_ net502 VPWR _1490_ VGND _1488_ _1489_ sg13g2_o21ai_1
X_5582_ _2297_ net1415 _2296_ VPWR VGND sg13g2_nand2_1
X_4533_ net385 VPWR _1434_ VGND net1477 net1532 sg13g2_o21ai_1
XFILLER_8_881 VPWR VGND sg13g2_decap_8
Xhold325 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[0\] VPWR VGND net1082
+ sg13g2_dlygate4sd3_1
Xhold314 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[8\] VPWR VGND net1071
+ sg13g2_dlygate4sd3_1
Xhold303 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[5\] VPWR VGND net1060
+ sg13g2_dlygate4sd3_1
Xhold336 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[0\] VPWR VGND net1093 sg13g2_dlygate4sd3_1
Xhold347 _1115_ VPWR VGND net1104 sg13g2_dlygate4sd3_1
Xhold369 _0336_ VPWR VGND net1126 sg13g2_dlygate4sd3_1
Xhold358 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[9\] VPWR VGND net1115
+ sg13g2_dlygate4sd3_1
X_6203_ net759 net426 _0441_ VPWR VGND sg13g2_nor2_1
X_4464_ net486 VPWR _1376_ VGND _1374_ _1375_ sg13g2_o21ai_1
X_4395_ _1315_ _1316_ _1317_ VPWR VGND sg13g2_nor2b_1
X_6134_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[3\] _2759_
+ _2760_ VPWR VGND sg13g2_and2_1
X_6065_ _2701_ net1318 _2699_ VPWR VGND sg13g2_xnor2_1
X_5016_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].y_shr\[10\] VPWR
+ _1835_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].z_sign _1833_
+ sg13g2_o21ai_1
X_6704__537 VPWR VGND net721 sg13g2_tiehi
X_5918_ VGND VPWR _2574_ net1249 _0393_ _2581_ sg13g2_a21oi_1
X_6898_ net733 VGND VPWR _0526_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[5\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_33_clk clknet_4_13_0_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
X_5849_ _2523_ net1346 _2521_ VPWR VGND sg13g2_xnor2_1
XFILLER_42_58 VPWR VGND sg13g2_fill_1
XFILLER_6_818 VPWR VGND sg13g2_decap_8
XFILLER_27_1023 VPWR VGND sg13g2_decap_4
XFILLER_18_947 VPWR VGND sg13g2_decap_8
XFILLER_45_799 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_24_clk clknet_4_7_0_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
XFILLER_5_884 VPWR VGND sg13g2_decap_8
X_4180_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[10\] VPWR _1138_ VGND
+ _1130_ _1131_ sg13g2_o21ai_1
X_6821_ net604 VGND VPWR net1299 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[1\]
+ clknet_leaf_62_clk sg13g2_dfrbpq_2
XFILLER_35_232 VPWR VGND sg13g2_fill_2
XFILLER_36_766 VPWR VGND sg13g2_fill_2
X_6752_ net673 VGND VPWR _0361_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[6\]
+ clknet_leaf_48_clk sg13g2_dfrbpq_2
X_3964_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[1\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt_sum\[5\]
+ _0965_ VPWR VGND sg13g2_xor2_1
Xclkbuf_leaf_15_clk clknet_4_4_0_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
X_3895_ _0914_ net1056 _0916_ VPWR VGND sg13g2_xor2_1
X_5703_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[10\] net412 _2394_
+ _2401_ VPWR VGND sg13g2_a21o_1
X_6683_ net756 VGND VPWR net1096 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[4\]
+ clknet_leaf_45_clk sg13g2_dfrbpq_1
X_5634_ _2342_ _2336_ net1194 VPWR VGND sg13g2_nand2b_1
X_6402__375 VPWR VGND net559 sg13g2_tiehi
X_5565_ _2282_ net1302 _2280_ VPWR VGND sg13g2_xnor2_1
Xhold100 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[0\] VPWR VGND net857 sg13g2_dlygate4sd3_1
X_4516_ _1419_ _1420_ _0152_ VPWR VGND sg13g2_nor2b_1
Xhold144 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[7\] VPWR VGND net901 sg13g2_dlygate4sd3_1
Xhold111 _0017_ VPWR VGND net868 sg13g2_dlygate4sd3_1
Xhold133 _0872_ VPWR VGND net890 sg13g2_dlygate4sd3_1
Xhold122 u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[0\] VPWR VGND net879 sg13g2_dlygate4sd3_1
X_5496_ net524 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[1\] _2226_
+ VPWR VGND sg13g2_nor2b_1
Xhold166 _1305_ VPWR VGND net923 sg13g2_dlygate4sd3_1
Xhold177 _2269_ VPWR VGND net934 sg13g2_dlygate4sd3_1
Xhold155 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[5\]\[0\] VPWR VGND net912
+ sg13g2_dlygate4sd3_1
X_4447_ _1357_ _1358_ _1361_ VPWR VGND sg13g2_nor2_1
Xhold188 _0016_ VPWR VGND net945 sg13g2_dlygate4sd3_1
Xhold199 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[8\] VPWR VGND net956
+ sg13g2_dlygate4sd3_1
X_6117_ _2745_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[3\] _2744_
+ VPWR VGND sg13g2_xnor2_1
X_4378_ VGND VPWR _1301_ _1302_ _0131_ _1303_ sg13g2_a21oi_1
X_6048_ net1209 _2685_ _2686_ VPWR VGND sg13g2_nor2_1
XFILLER_15_906 VPWR VGND sg13g2_decap_8
XFILLER_23_950 VPWR VGND sg13g2_decap_8
X_6854__378 VPWR VGND net562 sg13g2_tiehi
X_6518__204 VPWR VGND net204 sg13g2_tiehi
XFILLER_2_865 VPWR VGND sg13g2_decap_8
XFILLER_17_287 VPWR VGND sg13g2_fill_1
XFILLER_14_983 VPWR VGND sg13g2_decap_8
XFILLER_20_408 VPWR VGND sg13g2_fill_2
X_3680_ _0645_ _0703_ _0732_ _0733_ VPWR VGND sg13g2_nor3_1
X_5350_ _2101_ _2102_ _0304_ VPWR VGND sg13g2_nor2b_1
X_4301_ _0116_ net501 net1568 _1241_ VPWR VGND sg13g2_and3_1
X_5281_ net1473 net528 _2045_ VPWR VGND sg13g2_xor2_1
X_4232_ net382 VPWR _1182_ VGND net1300 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[5\]
+ sg13g2_o21ai_1
Xclkbuf_leaf_4_clk clknet_4_1_0_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_4163_ _0582_ VPWR _1123_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[6\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[7\] sg13g2_o21ai_1
X_4094_ net419 _1070_ _0079_ VPWR VGND sg13g2_nor2_1
X_6740__501 VPWR VGND net685 sg13g2_tiehi
X_4996_ _1814_ VPWR _1819_ VGND net1186 net398 sg13g2_o21ai_1
X_6804_ net621 VGND VPWR _0413_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].z_sign
+ clknet_leaf_9_clk sg13g2_dfrbpq_2
XFILLER_24_747 VPWR VGND sg13g2_fill_1
X_3947_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[10\] _0947_ _0948_
+ VPWR VGND sg13g2_nor2b_1
X_6735_ net690 VGND VPWR net1414 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[6\]
+ clknet_leaf_55_clk sg13g2_dfrbpq_1
XFILLER_17_1011 VPWR VGND sg13g2_decap_8
X_6666_ net56 VGND VPWR _0275_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[6\]\[0\]
+ clknet_leaf_51_clk sg13g2_dfrbpq_1
XFILLER_20_975 VPWR VGND sg13g2_decap_8
X_3878_ net419 net1094 _0031_ VPWR VGND sg13g2_nor2_1
X_5617_ net1335 _2327_ _0346_ VPWR VGND sg13g2_nor2b_1
X_6597_ net125 VGND VPWR _0206_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[8\]
+ clknet_leaf_26_clk sg13g2_dfrbpq_1
X_5548_ VGND VPWR _0553_ net811 _0337_ _2267_ sg13g2_a21oi_1
X_5479_ VGND VPWR _2213_ _2208_ _2205_ sg13g2_or2_1
Xfanout421 net422 net421 VPWR VGND sg13g2_buf_8
Xfanout432 net434 net432 VPWR VGND sg13g2_buf_8
Xfanout410 net411 net410 VPWR VGND sg13g2_buf_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
Xfanout443 net451 net443 VPWR VGND sg13g2_buf_8
Xfanout454 net456 net454 VPWR VGND sg13g2_buf_8
Xfanout465 net466 net465 VPWR VGND sg13g2_buf_8
XFILLER_19_508 VPWR VGND sg13g2_fill_1
Xfanout476 net491 net476 VPWR VGND sg13g2_buf_8
Xfanout487 net490 net487 VPWR VGND sg13g2_buf_1
Xfanout498 net500 net498 VPWR VGND sg13g2_buf_8
XFILLER_15_714 VPWR VGND sg13g2_fill_1
XFILLER_11_975 VPWR VGND sg13g2_decap_8
XFILLER_10_485 VPWR VGND sg13g2_fill_2
XFILLER_7_946 VPWR VGND sg13g2_decap_8
XFILLER_9_1009 VPWR VGND sg13g2_decap_8
XFILLER_1_183 VPWR VGND sg13g2_fill_1
XFILLER_38_839 VPWR VGND sg13g2_fill_1
XFILLER_18_552 VPWR VGND sg13g2_fill_1
X_4850_ _1689_ _1690_ _1694_ _1697_ VPWR VGND sg13g2_or3_1
X_3801_ _0636_ _0846_ _0011_ VPWR VGND sg13g2_nor2_1
X_4781_ net536 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[9\] _1639_
+ VPWR VGND sg13g2_nor2b_1
X_6520_ net202 VGND VPWR net1111 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[8\]
+ clknet_leaf_42_clk sg13g2_dfrbpq_1
X_3732_ _0785_ _0773_ _0784_ VPWR VGND sg13g2_nand2_1
X_6451_ net291 VGND VPWR net949 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[4\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_2
X_3663_ _0716_ _0704_ _0712_ VPWR VGND sg13g2_xnor2_1
X_6913__272 VPWR VGND net272 sg13g2_tiehi
X_6382_ VGND VPWR _2873_ _2877_ _0462_ _2878_ sg13g2_a21oi_1
X_5402_ _2132_ net1233 _2147_ VPWR VGND sg13g2_xor2_1
X_5333_ _2079_ VPWR _2087_ VGND net521 _0555_ sg13g2_o21ai_1
X_3594_ net546 u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[8\] u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[8\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[8\] net535 net544 _0647_
+ VPWR VGND sg13g2_mux4_1
X_5264_ _2034_ _0567_ _2007_ VPWR VGND sg13g2_xnor2_1
X_5195_ VGND VPWR _1968_ _1973_ _1975_ net439 sg13g2_a21oi_1
X_4215_ _1167_ _1168_ _0103_ VPWR VGND sg13g2_nor2b_1
X_4146_ _1108_ VPWR _1110_ VGND net533 _0591_ sg13g2_o21ai_1
X_6508__214 VPWR VGND net214 sg13g2_tiehi
X_4077_ _1058_ net849 _1060_ VPWR VGND sg13g2_xor2_1
X_4979_ _1805_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[7\] net397
+ VPWR VGND sg13g2_xnor2_1
X_6439__308 VPWR VGND net308 sg13g2_tiehi
Xclkload3 clknet_4_5_0_clk clkload3/X VPWR VGND sg13g2_buf_8
X_6718_ net707 VGND VPWR net853 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[1\]
+ clknet_leaf_32_clk sg13g2_dfrbpq_1
X_6649_ net73 VGND VPWR _0258_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[10\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_1
X_6515__207 VPWR VGND net207 sg13g2_tiehi
XFILLER_4_916 VPWR VGND sg13g2_decap_8
XFILLER_47_669 VPWR VGND sg13g2_fill_2
XFILLER_15_533 VPWR VGND sg13g2_fill_1
XFILLER_43_886 VPWR VGND sg13g2_fill_1
XFILLER_15_577 VPWR VGND sg13g2_decap_4
XFILLER_30_558 VPWR VGND sg13g2_fill_1
X_6730__511 VPWR VGND net695 sg13g2_tiehi
X_4000_ _0999_ net980 net376 VPWR VGND sg13g2_nand2_1
XFILLER_27_4 VPWR VGND sg13g2_fill_1
X_5951_ _2610_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[11\] _2609_
+ VPWR VGND sg13g2_xnor2_1
X_6839__402 VPWR VGND net586 sg13g2_tiehi
X_4902_ _1734_ VPWR _1740_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[7\]
+ net389 sg13g2_o21ai_1
X_5882_ VGND VPWR _2545_ _2549_ _2551_ _2548_ sg13g2_a21oi_1
X_6874__337 VPWR VGND net337 sg13g2_tiehi
XFILLER_21_525 VPWR VGND sg13g2_fill_1
X_4833_ net426 _1682_ _1683_ _0206_ VPWR VGND sg13g2_nor3_1
X_4764_ _1625_ net401 _1514_ VPWR VGND sg13g2_nand2b_1
XFILLER_14_1025 VPWR VGND sg13g2_decap_4
X_3715_ _0768_ _0766_ _0767_ VPWR VGND sg13g2_xnor2_1
X_6503_ net219 VGND VPWR _0112_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[4\]
+ clknet_leaf_45_clk sg13g2_dfrbpq_1
X_4695_ _1567_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[1\] _1565_
+ VPWR VGND sg13g2_xnor2_1
X_6434_ net313 VGND VPWR _0043_ u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[0\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
X_3646_ net407 net409 _0699_ VPWR VGND sg13g2_xor2_1
X_3577_ _0634_ net878 net859 VPWR VGND sg13g2_nand2b_1
X_6365_ net958 _2917_ _2920_ VPWR VGND sg13g2_nor2_1
X_6296_ _2883_ _2889_ _2870_ _2891_ VPWR VGND sg13g2_nand3_1
X_5316_ net971 _2071_ _0300_ VPWR VGND sg13g2_nor2b_1
X_5247_ _2020_ _2014_ _2017_ VPWR VGND sg13g2_nand2_1
Xhold15 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[0\] VPWR VGND net772
+ sg13g2_dlygate4sd3_1
Xhold26 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[3\] VPWR VGND net783
+ sg13g2_dlygate4sd3_1
Xhold37 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[9\] VPWR VGND net794
+ sg13g2_dlygate4sd3_1
Xhold48 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[4\] VPWR VGND net805
+ sg13g2_dlygate4sd3_1
Xhold59 _0488_ VPWR VGND net816 sg13g2_dlygate4sd3_1
X_5178_ VGND VPWR _1958_ _1959_ _0274_ _1960_ sg13g2_a21oi_1
XFILLER_28_113 VPWR VGND sg13g2_fill_1
X_4129_ _1094_ _1095_ _1096_ VPWR VGND sg13g2_nor2_1
XFILLER_25_853 VPWR VGND sg13g2_fill_2
XFILLER_4_713 VPWR VGND sg13g2_decap_8
XFILLER_3_256 VPWR VGND sg13g2_fill_2
XFILLER_0_941 VPWR VGND sg13g2_decap_8
XFILLER_48_934 VPWR VGND sg13g2_fill_2
X_6628__94 VPWR VGND net94 sg13g2_tiehi
XFILLER_16_886 VPWR VGND sg13g2_decap_8
XFILLER_37_1003 VPWR VGND sg13g2_fill_1
X_3500_ VPWR _0570_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[9\] VGND
+ sg13g2_inv_1
Xhold507 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[2\] VPWR VGND net1264
+ sg13g2_dlygate4sd3_1
Xhold518 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[4\] VPWR VGND net1275
+ sg13g2_dlygate4sd3_1
X_4480_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[2\] _1388_ _1389_
+ VPWR VGND sg13g2_and2_1
Xhold529 _0325_ VPWR VGND net1286 sg13g2_dlygate4sd3_1
X_6150_ net1420 _2773_ _2774_ VPWR VGND sg13g2_and2_1
X_5101_ _1892_ _1893_ _1894_ VPWR VGND sg13g2_nor2b_1
X_6081_ _2715_ _0623_ _2713_ VPWR VGND sg13g2_xnor2_1
X_5032_ _1847_ _1848_ _1844_ _1849_ VPWR VGND sg13g2_nand3_1
X_6505__217 VPWR VGND net217 sg13g2_tiehi
XFILLER_25_138 VPWR VGND sg13g2_fill_1
X_5934_ net425 _2594_ _2595_ _0395_ VPWR VGND sg13g2_nor3_1
X_5865_ _2537_ net1326 _2535_ VPWR VGND sg13g2_xnor2_1
X_4816_ _1668_ VPWR _1669_ VGND _1664_ _1665_ sg13g2_o21ai_1
X_5796_ _2476_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[1\]
+ _2475_ VPWR VGND sg13g2_xnor2_1
X_4747_ _1610_ _1611_ _0192_ VPWR VGND sg13g2_nor2_1
XFILLER_31_27 VPWR VGND sg13g2_fill_2
X_4678_ VGND VPWR u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[2\]
+ net394 _1553_ _1552_ sg13g2_a21oi_1
X_6417_ net346 VGND VPWR net1032 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[6\] clknet_leaf_66_clk
+ sg13g2_dfrbpq_2
X_3629_ VGND VPWR net405 _0647_ _0682_ _0642_ sg13g2_a21oi_1
X_6348_ _0547_ _2906_ _2909_ VPWR VGND sg13g2_and2_1
XFILLER_1_749 VPWR VGND sg13g2_decap_8
XFILLER_49_709 VPWR VGND sg13g2_fill_1
X_6279_ VGND VPWR net939 net1070 _2879_ _2864_ sg13g2_a21oi_1
XFILLER_17_639 VPWR VGND sg13g2_fill_2
X_6720__521 VPWR VGND net705 sg13g2_tiehi
X_6625__97 VPWR VGND net97 sg13g2_tiehi
XFILLER_21_60 VPWR VGND sg13g2_fill_2
X_6829__412 VPWR VGND net596 sg13g2_tiehi
XFILLER_36_948 VPWR VGND sg13g2_fill_2
X_3980_ _0981_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[15\] _0980_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_16_683 VPWR VGND sg13g2_fill_2
X_6836__405 VPWR VGND net589 sg13g2_tiehi
X_5650_ net474 VPWR _2355_ VGND _2349_ _2354_ sg13g2_o21ai_1
XFILLER_15_193 VPWR VGND sg13g2_fill_2
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
X_4601_ net832 net540 _1489_ VPWR VGND sg13g2_xor2_1
X_5581_ _2294_ _2295_ _2296_ VPWR VGND sg13g2_nor2b_1
X_4532_ _1433_ _1428_ _1430_ VPWR VGND sg13g2_nand2_1
XFILLER_8_860 VPWR VGND sg13g2_decap_8
XFILLER_7_51 VPWR VGND sg13g2_fill_2
XFILLER_11_1017 VPWR VGND sg13g2_decap_8
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
Xhold326 _1638_ VPWR VGND net1083 sg13g2_dlygate4sd3_1
Xhold315 _2848_ VPWR VGND net1072 sg13g2_dlygate4sd3_1
Xhold304 _0088_ VPWR VGND net1061 sg13g2_dlygate4sd3_1
X_4463_ _1375_ net1287 net387 VPWR VGND sg13g2_xnor2_1
Xhold337 _0903_ VPWR VGND net1094 sg13g2_dlygate4sd3_1
Xhold348 _0096_ VPWR VGND net1105 sg13g2_dlygate4sd3_1
Xhold359 _0092_ VPWR VGND net1116 sg13g2_dlygate4sd3_1
X_6202_ net466 net761 _0440_ VPWR VGND sg13g2_and2_1
X_4394_ _1313_ _1314_ _0604_ _1316_ VPWR VGND sg13g2_nand3_1
X_6133_ _2759_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[5\] _2758_
+ VPWR VGND sg13g2_xnor2_1
X_6064_ _2700_ net1318 _2699_ VPWR VGND sg13g2_nand2_1
X_5015_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].z_sign u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].y_shr\[10\]
+ _1833_ _1834_ VPWR VGND sg13g2_nor3_1
XFILLER_42_907 VPWR VGND sg13g2_fill_2
X_5917_ net457 VPWR _2581_ VGND _2574_ _2580_ sg13g2_o21ai_1
X_6897_ net732 VGND VPWR _0525_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[4\]
+ clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5848_ _2522_ net1346 _2521_ VPWR VGND sg13g2_nand2_1
XFILLER_10_859 VPWR VGND sg13g2_decap_8
X_5779_ VGND VPWR _2460_ _2462_ _2464_ net425 sg13g2_a21oi_1
XFILLER_27_1002 VPWR VGND sg13g2_decap_8
XFILLER_18_926 VPWR VGND sg13g2_decap_8
XFILLER_44_299 VPWR VGND sg13g2_fill_1
XFILLER_44_266 VPWR VGND sg13g2_fill_1
XFILLER_32_439 VPWR VGND sg13g2_fill_2
XFILLER_41_973 VPWR VGND sg13g2_fill_1
XFILLER_5_863 VPWR VGND sg13g2_decap_8
X_6820_ net605 VGND VPWR _0429_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[0\]
+ clknet_leaf_62_clk sg13g2_dfrbpq_2
X_6751_ net674 VGND VPWR net1451 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[5\]
+ clknet_leaf_57_clk sg13g2_dfrbpq_1
X_3963_ _0964_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[3\] _0942_
+ VPWR VGND sg13g2_xnor2_1
X_3894_ net420 net1004 _0915_ _0035_ VPWR VGND sg13g2_nor3_1
X_5702_ _2396_ VPWR _2400_ VGND _2393_ _2398_ sg13g2_o21ai_1
X_6682_ net40 VGND VPWR _0291_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[3\]
+ clknet_leaf_45_clk sg13g2_dfrbpq_1
X_5633_ _2338_ _2334_ _2337_ _2341_ VPWR VGND sg13g2_a21o_1
X_5564_ _2281_ net1302 _2280_ VPWR VGND sg13g2_nand2_1
X_4515_ VGND VPWR _1415_ _1418_ _1420_ net438 sg13g2_a21oi_1
Xhold101 _0020_ VPWR VGND net858 sg13g2_dlygate4sd3_1
Xhold112 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[7\] VPWR VGND net869 sg13g2_dlygate4sd3_1
Xhold134 _0019_ VPWR VGND net891 sg13g2_dlygate4sd3_1
Xhold123 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[10\] VPWR VGND net880
+ sg13g2_dlygate4sd3_1
X_5495_ net852 net432 _0326_ VPWR VGND sg13g2_nor2_1
Xhold167 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[1\] VPWR VGND
+ net924 sg13g2_dlygate4sd3_1
X_6710__531 VPWR VGND net715 sg13g2_tiehi
Xhold156 _1962_ VPWR VGND net913 sg13g2_dlygate4sd3_1
Xhold145 _0038_ VPWR VGND net902 sg13g2_dlygate4sd3_1
X_4446_ VGND VPWR _1358_ _1359_ _0142_ _1360_ sg13g2_a21oi_1
Xhold189 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[0\] VPWR VGND net946
+ sg13g2_dlygate4sd3_1
Xhold178 _0338_ VPWR VGND net935 sg13g2_dlygate4sd3_1
X_4377_ net501 VPWR _1303_ VGND _1301_ _1302_ sg13g2_o21ai_1
X_6116_ net507 _2743_ _2744_ VPWR VGND sg13g2_nor2_1
X_6923__252 VPWR VGND net252 sg13g2_tiehi
X_6047_ _2684_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[5\]
+ _2685_ VPWR VGND sg13g2_xor2_1
XFILLER_2_1026 VPWR VGND sg13g2_fill_2
XFILLER_26_222 VPWR VGND sg13g2_fill_2
XFILLER_42_737 VPWR VGND sg13g2_fill_2
X_6819__422 VPWR VGND net606 sg13g2_tiehi
XFILLER_41_269 VPWR VGND sg13g2_fill_1
XFILLER_10_667 VPWR VGND sg13g2_fill_1
Xhold690 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[3\] VPWR VGND net1447
+ sg13g2_dlygate4sd3_1
XFILLER_2_844 VPWR VGND sg13g2_decap_8
X_6826__415 VPWR VGND net599 sg13g2_tiehi
XFILLER_49_369 VPWR VGND sg13g2_fill_2
XFILLER_17_222 VPWR VGND sg13g2_fill_1
XFILLER_17_277 VPWR VGND sg13g2_fill_1
XFILLER_33_748 VPWR VGND sg13g2_fill_2
XFILLER_14_962 VPWR VGND sg13g2_decap_8
X_6833__408 VPWR VGND net592 sg13g2_tiehi
XFILLER_9_421 VPWR VGND sg13g2_fill_2
X_4300_ _1239_ VPWR _1241_ VGND _1235_ _1238_ sg13g2_o21ai_1
X_5280_ _2044_ net415 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[5\]
+ VPWR VGND sg13g2_nand2_1
X_4231_ _1172_ _1173_ _1178_ _1181_ VPWR VGND sg13g2_nor3_1
X_4162_ _1119_ VPWR _1122_ VGND _1115_ _1120_ sg13g2_o21ai_1
X_4093_ _1070_ net865 _1069_ VPWR VGND sg13g2_xnor2_1
X_6803_ net622 VGND VPWR _0412_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[10\]
+ clknet_leaf_9_clk sg13g2_dfrbpq_1
X_4995_ _1818_ net1052 net399 VPWR VGND sg13g2_xnor2_1
X_6734_ net691 VGND VPWR net1416 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[5\]
+ clknet_leaf_55_clk sg13g2_dfrbpq_2
X_3946_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[8\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[9\]
+ _0946_ _0947_ VPWR VGND sg13g2_nor3_1
X_3877_ _0902_ VPWR _0903_ VGND net1093 _0901_ sg13g2_o21ai_1
XFILLER_20_954 VPWR VGND sg13g2_decap_8
X_6665_ net57 VGND VPWR net1409 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[12\]
+ clknet_leaf_50_clk sg13g2_dfrbpq_2
X_5616_ VGND VPWR _2320_ _2325_ _2327_ net431 sg13g2_a21oi_1
X_6596_ net126 VGND VPWR net1092 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[7\]
+ clknet_leaf_28_clk sg13g2_dfrbpq_2
X_5547_ VGND VPWR net1125 _2266_ _0336_ _2267_ sg13g2_a21oi_1
X_5478_ _2206_ net1483 _2212_ VPWR VGND sg13g2_xor2_1
X_6884__317 VPWR VGND net317 sg13g2_tiehi
X_4429_ _1340_ _1338_ _1344_ _1347_ VPWR VGND sg13g2_a21o_1
Xfanout400 net401 net400 VPWR VGND sg13g2_buf_8
XFILLER_48_14 VPWR VGND sg13g2_decap_8
Xfanout422 net423 net422 VPWR VGND sg13g2_buf_8
Xfanout411 _0600_ net411 VPWR VGND sg13g2_buf_8
Xfanout444 net447 net444 VPWR VGND sg13g2_buf_8
Xfanout455 net456 net455 VPWR VGND sg13g2_buf_1
XFILLER_24_1016 VPWR VGND sg13g2_decap_8
XFILLER_24_1027 VPWR VGND sg13g2_fill_2
Xfanout433 net434 net433 VPWR VGND sg13g2_buf_8
Xfanout466 net473 net466 VPWR VGND sg13g2_buf_8
Xfanout488 net490 net488 VPWR VGND sg13g2_buf_8
Xfanout477 net478 net477 VPWR VGND sg13g2_buf_8
X_6682__40 VPWR VGND net40 sg13g2_tiehi
Xfanout499 net500 net499 VPWR VGND sg13g2_buf_1
XFILLER_42_523 VPWR VGND sg13g2_fill_1
XFILLER_30_718 VPWR VGND sg13g2_fill_1
XFILLER_7_925 VPWR VGND sg13g2_decap_8
XFILLER_11_954 VPWR VGND sg13g2_decap_8
XFILLER_6_413 VPWR VGND sg13g2_fill_1
XFILLER_29_8 VPWR VGND sg13g2_fill_1
X_4780_ net432 net1083 _0198_ VPWR VGND sg13g2_nor2_2
X_3800_ net451 VPWR _0846_ VGND _0651_ _0685_ sg13g2_o21ai_1
X_3731_ _0784_ _0750_ _0782_ VPWR VGND sg13g2_xnor2_1
X_6450_ net293 VGND VPWR net955 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[3\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_2
X_3662_ _0713_ _0714_ _0715_ VPWR VGND sg13g2_nor2_1
Xclkload10 clknet_4_13_0_clk clkload10/X VPWR VGND sg13g2_buf_8
X_6381_ VGND VPWR _2860_ _2862_ _0457_ net421 sg13g2_a21oi_1
X_5401_ _2143_ VPWR _2146_ VGND _2141_ _2142_ sg13g2_o21ai_1
X_3593_ net546 u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[9\] u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[9\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[9\] net535 net544 _0646_
+ VPWR VGND sg13g2_mux4_1
X_5332_ VGND VPWR _2078_ _2082_ _2086_ _2081_ sg13g2_a21oi_1
XFILLER_47_1027 VPWR VGND sg13g2_fill_2
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_6809__432 VPWR VGND net616 sg13g2_tiehi
X_5263_ _2031_ _2032_ _2025_ _2033_ VPWR VGND sg13g2_nand3_1
X_5194_ _1968_ _1973_ _1974_ VPWR VGND sg13g2_nor2_1
X_4214_ VGND VPWR _1165_ _1166_ _1168_ net433 sg13g2_a21oi_1
XFILLER_28_306 VPWR VGND sg13g2_fill_2
X_4145_ VGND VPWR _1106_ _1107_ _0092_ _1109_ sg13g2_a21oi_1
X_4076_ net849 net919 _1054_ _1059_ VPWR VGND sg13g2_nor3_1
XFILLER_24_512 VPWR VGND sg13g2_fill_1
XFILLER_11_217 VPWR VGND sg13g2_fill_1
X_6816__425 VPWR VGND net609 sg13g2_tiehi
X_4978_ VGND VPWR net1122 net397 _1804_ _1802_ sg13g2_a21oi_1
X_6717_ net708 VGND VPWR _0326_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[0\]
+ clknet_leaf_35_clk sg13g2_dfrbpq_1
Xclkload4 clknet_4_6_0_clk clkload4/X VPWR VGND sg13g2_buf_8
X_3929_ net982 net1012 _0532_ _0931_ VPWR VGND net918 sg13g2_nand4_1
X_6648_ net74 VGND VPWR _0257_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[9\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_1
XFILLER_30_1020 VPWR VGND sg13g2_decap_8
X_6579_ net143 VGND VPWR _0188_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[4\]
+ clknet_leaf_34_clk sg13g2_dfrbpq_2
XFILLER_3_427 VPWR VGND sg13g2_fill_1
XFILLER_8_1021 VPWR VGND sg13g2_decap_8
X_6823__418 VPWR VGND net602 sg13g2_tiehi
XFILLER_7_799 VPWR VGND sg13g2_decap_8
XFILLER_3_983 VPWR VGND sg13g2_decap_8
X_5950_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[10\] net414 _2603_
+ _2609_ VPWR VGND sg13g2_a21o_1
XFILLER_37_169 VPWR VGND sg13g2_fill_2
X_4901_ VGND VPWR _1737_ _1738_ _0218_ _1739_ sg13g2_a21oi_1
XFILLER_34_843 VPWR VGND sg13g2_fill_1
X_5881_ VGND VPWR _2545_ _2549_ _0387_ _2550_ sg13g2_a21oi_1
X_4832_ _1681_ _1680_ _1683_ VPWR VGND sg13g2_nor2b_1
X_4763_ _1624_ _1615_ _1622_ VPWR VGND sg13g2_nand2_1
XFILLER_14_1004 VPWR VGND sg13g2_decap_8
X_3714_ VGND VPWR _0679_ _0696_ _0767_ _0745_ sg13g2_a21oi_1
X_4694_ _1566_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[1\] _1565_
+ VPWR VGND sg13g2_nand2_1
X_6502_ net220 VGND VPWR _0111_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[3\]
+ clknet_leaf_32_clk sg13g2_dfrbpq_1
X_6433_ net314 VGND VPWR _0042_ u_angle_cordic_12b_pmod.u_vga_top.pixel_clk_en clknet_leaf_65_clk
+ sg13g2_dfrbpq_2
X_3645_ _0698_ _0679_ _0696_ VPWR VGND sg13g2_xnor2_1
X_3576_ _0633_ net442 net822 VPWR VGND sg13g2_nand2_1
X_6364_ net958 _2917_ _2919_ VPWR VGND sg13g2_and2_1
X_6295_ _2888_ _2890_ _0470_ VPWR VGND sg13g2_nor2_1
X_5315_ net477 VPWR _2072_ VGND net970 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[0\]
+ sg13g2_o21ai_1
X_5246_ net379 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[4\]
+ _2019_ VPWR VGND sg13g2_xor2_1
Xhold27 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[3\] VPWR VGND net784
+ sg13g2_dlygate4sd3_1
Xhold38 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[10\] VPWR VGND net795
+ sg13g2_dlygate4sd3_1
XFILLER_29_38 VPWR VGND sg13g2_fill_1
Xhold16 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[4\] VPWR VGND net773
+ sg13g2_dlygate4sd3_1
Xhold49 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[0\] VPWR VGND net806
+ sg13g2_dlygate4sd3_1
X_5177_ net492 VPWR _1960_ VGND _1958_ _1959_ sg13g2_o21ai_1
X_6445__302 VPWR VGND net302 sg13g2_tiehi
XFILLER_28_147 VPWR VGND sg13g2_fill_1
X_4128_ _1087_ VPWR _1095_ VGND net533 _0589_ sg13g2_o21ai_1
X_4059_ _0532_ net423 _0082_ VPWR VGND sg13g2_nor2_1
X_6521__201 VPWR VGND net201 sg13g2_tiehi
XFILLER_36_191 VPWR VGND sg13g2_fill_2
XFILLER_8_508 VPWR VGND sg13g2_fill_1
XFILLER_12_548 VPWR VGND sg13g2_fill_2
XFILLER_4_769 VPWR VGND sg13g2_decap_8
XFILLER_0_920 VPWR VGND sg13g2_decap_8
XFILLER_0_997 VPWR VGND sg13g2_decap_8
XFILLER_19_125 VPWR VGND sg13g2_fill_1
XFILLER_34_117 VPWR VGND sg13g2_fill_1
XFILLER_30_389 VPWR VGND sg13g2_fill_2
XFILLER_11_592 VPWR VGND sg13g2_fill_2
XFILLER_7_563 VPWR VGND sg13g2_fill_1
Xhold508 _2738_ VPWR VGND net1265 sg13g2_dlygate4sd3_1
Xhold519 _0267_ VPWR VGND net1276 sg13g2_dlygate4sd3_1
X_6080_ _2714_ net1371 _2713_ VPWR VGND sg13g2_nand2b_1
XFILLER_3_780 VPWR VGND sg13g2_decap_8
X_5100_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[2\] _1891_
+ net415 _1893_ VPWR VGND sg13g2_nand3_1
X_5031_ _1848_ _0618_ _1842_ VPWR VGND sg13g2_xnor2_1
X_6806__435 VPWR VGND net619 sg13g2_tiehi
X_5933_ _2589_ _2593_ _2595_ VPWR VGND sg13g2_and2_1
X_5864_ _2535_ net1326 _2536_ VPWR VGND sg13g2_nor2b_1
X_4815_ net391 VPWR _1668_ VGND net1237 net1545 sg13g2_o21ai_1
X_5795_ net512 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[0\]
+ _2475_ VPWR VGND sg13g2_nor2b_1
X_4746_ _1611_ net489 net1459 VPWR VGND sg13g2_nand2_1
X_6813__428 VPWR VGND net612 sg13g2_tiehi
X_4677_ net432 _1551_ net1535 _0181_ VPWR VGND sg13g2_nor3_1
X_6416_ net348 VGND VPWR _0025_ u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[5\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_2
X_3628_ _0681_ net405 _0655_ VPWR VGND sg13g2_nand2_1
X_6347_ _0547_ _2906_ _2908_ VPWR VGND sg13g2_nor2_1
Xoutput17 net17 uio_out[7] VPWR VGND sg13g2_buf_1
XFILLER_1_728 VPWR VGND sg13g2_decap_8
X_3559_ net849 net451 _0524_ VPWR VGND sg13g2_and2_1
X_6278_ VGND VPWR _2873_ _2877_ _0459_ _2878_ sg13g2_a21oi_1
X_6412__356 VPWR VGND net356 sg13g2_tiehi
X_5229_ _2003_ _2004_ _0281_ VPWR VGND sg13g2_nor2_1
XFILLER_5_1024 VPWR VGND sg13g2_decap_4
XFILLER_45_938 VPWR VGND sg13g2_fill_2
XFILLER_0_794 VPWR VGND sg13g2_decap_8
XFILLER_31_676 VPWR VGND sg13g2_fill_1
X_4600_ VGND VPWR _0608_ net1185 _1488_ _1487_ sg13g2_a21oi_1
X_5580_ _0595_ VPWR _2295_ VGND net515 _2286_ sg13g2_o21ai_1
X_4531_ VGND VPWR _1430_ _1431_ _0155_ _1432_ sg13g2_a21oi_1
Xhold305 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[5\]\[1\] VPWR VGND net1062
+ sg13g2_dlygate4sd3_1
XFILLER_7_371 VPWR VGND sg13g2_fill_1
Xhold316 _0449_ VPWR VGND net1073 sg13g2_dlygate4sd3_1
X_4462_ VGND VPWR _1361_ _1371_ _1374_ _1373_ sg13g2_a21oi_1
X_6435__312 VPWR VGND net312 sg13g2_tiehi
X_6201_ VGND VPWR _2815_ net1282 _0439_ _2818_ sg13g2_a21oi_1
Xhold349 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[6\] VPWR VGND net1106
+ sg13g2_dlygate4sd3_1
Xhold327 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[5\] VPWR VGND net1084
+ sg13g2_dlygate4sd3_1
Xhold338 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[4\] VPWR VGND net1095
+ sg13g2_dlygate4sd3_1
X_6511__211 VPWR VGND net211 sg13g2_tiehi
X_4393_ VGND VPWR _1313_ _1314_ _1315_ _0604_ sg13g2_a21oi_1
X_6132_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[4\] net416 _2752_
+ _2758_ VPWR VGND sg13g2_a21o_1
X_6063_ _2699_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[7\]
+ _2698_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_220 VPWR VGND sg13g2_fill_2
X_5014_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].y_shr\[0\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].y_shr\[1\]
+ _1833_ VPWR VGND sg13g2_nor2_1
X_6442__305 VPWR VGND net305 sg13g2_tiehi
X_5916_ _2580_ net1248 _2577_ VPWR VGND sg13g2_xnor2_1
X_6893__544 VPWR VGND net728 sg13g2_tiehi
XFILLER_35_982 VPWR VGND sg13g2_fill_2
X_6896_ net731 VGND VPWR net850 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[3\]
+ clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5847_ _2520_ net1571 _2521_ VPWR VGND sg13g2_xor2_1
X_5778_ _2460_ _2462_ _2463_ VPWR VGND sg13g2_nor2_1
X_4729_ net1495 net400 _1596_ VPWR VGND sg13g2_and2_1
XFILLER_18_905 VPWR VGND sg13g2_decap_8
XFILLER_45_779 VPWR VGND sg13g2_fill_2
XFILLER_26_993 VPWR VGND sg13g2_decap_8
XFILLER_5_842 VPWR VGND sg13g2_decap_8
XFILLER_48_573 VPWR VGND sg13g2_fill_2
X_6803__438 VPWR VGND net622 sg13g2_tiehi
X_6750_ net675 VGND VPWR net1521 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[4\]
+ clknet_leaf_57_clk sg13g2_dfrbpq_2
XFILLER_44_790 VPWR VGND sg13g2_fill_1
X_5701_ VGND VPWR _2393_ _2398_ _0358_ _2399_ sg13g2_a21oi_1
X_3962_ _0944_ _0962_ _0963_ VPWR VGND sg13g2_nor2b_1
X_3893_ VPWR _0915_ _0914_ VGND sg13g2_inv_1
X_6681_ net41 VGND VPWR _0290_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[2\]
+ clknet_leaf_45_clk sg13g2_dfrbpq_1
X_5632_ net1468 _2340_ _0348_ VPWR VGND sg13g2_nor2b_1
X_5563_ _2280_ _0594_ _2279_ VPWR VGND sg13g2_xnor2_1
X_4514_ _1415_ _1418_ _1419_ VPWR VGND sg13g2_nor2_1
Xhold102 u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[10\] VPWR VGND net859 sg13g2_dlygate4sd3_1
Xhold113 _0868_ VPWR VGND net870 sg13g2_dlygate4sd3_1
Xhold135 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[2\] VPWR VGND net892 sg13g2_dlygate4sd3_1
X_5494_ VGND VPWR _2223_ _2224_ _0325_ _2225_ sg13g2_a21oi_1
Xhold124 _2914_ VPWR VGND net881 sg13g2_dlygate4sd3_1
Xhold168 _0057_ VPWR VGND net925 sg13g2_dlygate4sd3_1
Xhold157 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[8\] VPWR VGND net914 sg13g2_dlygate4sd3_1
Xhold146 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[10\] VPWR
+ VGND net903 sg13g2_dlygate4sd3_1
X_4445_ net486 VPWR _1360_ VGND _1358_ _1359_ sg13g2_o21ai_1
Xhold179 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[3\] VPWR VGND net936 sg13g2_dlygate4sd3_1
X_4376_ net818 net541 _1302_ VPWR VGND sg13g2_xor2_1
X_6115_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[1\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[2\]
+ _2743_ VPWR VGND sg13g2_nor2_1
X_6046_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[4\] net416
+ _2677_ _2684_ VPWR VGND sg13g2_a21o_1
XFILLER_2_1005 VPWR VGND sg13g2_decap_8
XFILLER_14_418 VPWR VGND sg13g2_fill_2
XFILLER_26_256 VPWR VGND sg13g2_fill_2
XFILLER_10_602 VPWR VGND sg13g2_fill_1
X_6879_ net327 VGND VPWR net816 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].z_sign
+ clknet_leaf_3_clk sg13g2_dfrbpq_1
XFILLER_23_985 VPWR VGND sg13g2_decap_8
XFILLER_2_823 VPWR VGND sg13g2_decap_8
Xhold680 _0397_ VPWR VGND net1437 sg13g2_dlygate4sd3_1
Xhold691 _0214_ VPWR VGND net1448 sg13g2_dlygate4sd3_1
XFILLER_14_941 VPWR VGND sg13g2_decap_8
X_6501__221 VPWR VGND net221 sg13g2_tiehi
X_4230_ VGND VPWR _1178_ _1179_ _0106_ _1180_ sg13g2_a21oi_1
X_4161_ VGND VPWR net1104 _1120_ _0096_ _1121_ sg13g2_a21oi_1
X_4092_ net420 _1068_ _1069_ _0078_ VPWR VGND sg13g2_nor3_1
X_6802_ net623 VGND VPWR net1155 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[9\]
+ clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_23_237 VPWR VGND sg13g2_fill_1
X_4994_ VGND VPWR _1814_ _1816_ _0233_ _1817_ sg13g2_a21oi_1
X_6733_ net692 VGND VPWR _0342_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[4\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_2
XFILLER_32_760 VPWR VGND sg13g2_fill_2
X_3945_ _0946_ _0945_ VPWR VGND u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[7\]
+ sg13g2_nand2b_2
XFILLER_20_933 VPWR VGND sg13g2_decap_8
X_6664_ net58 VGND VPWR net1292 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[11\]
+ clknet_leaf_49_clk sg13g2_dfrbpq_2
X_5615_ _2320_ _2325_ _2326_ VPWR VGND sg13g2_nor2_1
X_3876_ _0902_ net1093 _0884_ VPWR VGND sg13g2_nand2_1
X_6617__105 VPWR VGND net105 sg13g2_tiehi
X_6595_ net127 VGND VPWR _0204_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[6\]
+ clknet_leaf_29_clk sg13g2_dfrbpq_2
X_5546_ net479 VPWR _2267_ VGND net1125 _2266_ sg13g2_o21ai_1
X_5477_ _2211_ net1483 _2207_ VPWR VGND sg13g2_nand2_1
X_4428_ VGND VPWR _1338_ _1340_ _1346_ _1344_ sg13g2_a21oi_1
Xfanout401 _1592_ net401 VPWR VGND sg13g2_buf_8
Xfanout423 net440 net423 VPWR VGND sg13g2_buf_8
Xfanout412 _0592_ net412 VPWR VGND sg13g2_buf_8
Xfanout456 net473 net456 VPWR VGND sg13g2_buf_2
Xfanout434 net440 net434 VPWR VGND sg13g2_buf_8
Xfanout445 net447 net445 VPWR VGND sg13g2_buf_8
X_4359_ _1288_ _1283_ _1285_ _1287_ VPWR VGND sg13g2_and3_1
Xfanout489 net490 net489 VPWR VGND sg13g2_buf_1
Xfanout478 net480 net478 VPWR VGND sg13g2_buf_8
Xfanout467 net468 net467 VPWR VGND sg13g2_buf_8
X_6029_ net507 _2668_ _2669_ VPWR VGND sg13g2_nor2_1
X_6899__550 VPWR VGND net734 sg13g2_tiehi
XFILLER_11_933 VPWR VGND sg13g2_decap_8
XFILLER_7_904 VPWR VGND sg13g2_decap_8
XFILLER_2_697 VPWR VGND sg13g2_decap_8
X_3730_ _0750_ _0782_ _0783_ VPWR VGND sg13g2_nor2b_1
X_3661_ _0678_ _0661_ _0714_ VPWR VGND sg13g2_xor2_1
X_6380_ VGND VPWR _2860_ _2862_ _0456_ net421 sg13g2_a21oi_1
X_5400_ VGND VPWR _2141_ _2144_ _0311_ _2145_ sg13g2_a21oi_1
X_3592_ net407 net406 _0645_ VPWR VGND sg13g2_nor2_1
Xclkload11 clknet_4_14_0_clk clkload11/X VPWR VGND sg13g2_buf_8
X_5331_ net429 _2084_ _2085_ _0302_ VPWR VGND sg13g2_nor3_1
X_5262_ net379 VPWR _2032_ VGND net1227 net1314 sg13g2_o21ai_1
X_5193_ _1973_ net1337 _1971_ VPWR VGND sg13g2_xnor2_1
X_4213_ _1165_ _1166_ _1167_ VPWR VGND sg13g2_nor2_1
X_4144_ _1109_ net501 _1108_ VPWR VGND sg13g2_nand2_1
XFILLER_29_808 VPWR VGND sg13g2_fill_1
X_4075_ net919 _1054_ _1058_ VPWR VGND sg13g2_nor2_1
X_6716_ net709 VGND VPWR net1286 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[10\]
+ clknet_leaf_49_clk sg13g2_dfrbpq_1
X_4977_ _1802_ _1803_ _0230_ VPWR VGND sg13g2_nor2b_1
Xclkload5 clknet_4_7_0_clk clkload5/X VPWR VGND sg13g2_buf_8
X_3928_ net952 VPWR _0930_ VGND net961 _0929_ sg13g2_o21ai_1
X_3859_ _0888_ net1031 _0026_ VPWR VGND sg13g2_nor2_1
X_6647_ net75 VGND VPWR _0256_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[8\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
X_6578_ net144 VGND VPWR net1312 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[3\]
+ clknet_leaf_35_clk sg13g2_dfrbpq_1
X_5529_ _2253_ net523 net1156 VPWR VGND sg13g2_xnor2_1
XFILLER_8_1000 VPWR VGND sg13g2_decap_8
XFILLER_27_362 VPWR VGND sg13g2_fill_2
X_6422__336 VPWR VGND net336 sg13g2_tiehi
XFILLER_7_767 VPWR VGND sg13g2_decap_4
XFILLER_6_211 VPWR VGND sg13g2_fill_1
XFILLER_3_962 VPWR VGND sg13g2_decap_8
XFILLER_41_8 VPWR VGND sg13g2_fill_1
X_6607__115 VPWR VGND net115 sg13g2_tiehi
X_6466__263 VPWR VGND net263 sg13g2_tiehi
X_4900_ net485 VPWR _1739_ VGND _1737_ _1738_ sg13g2_o21ai_1
X_5880_ net459 VPWR _2550_ VGND _2545_ _2549_ sg13g2_o21ai_1
X_4831_ net1516 _1681_ _1682_ VPWR VGND sg13g2_nor2b_1
X_4762_ VGND VPWR _1621_ _1622_ _0195_ _1623_ sg13g2_a21oi_1
X_3713_ _0763_ _0748_ _0766_ VPWR VGND sg13g2_xor2_1
X_6501_ net221 VGND VPWR _0110_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[2\]
+ clknet_leaf_46_clk sg13g2_dfrbpq_1
X_4693_ _1565_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[1\]
+ _1564_ VPWR VGND sg13g2_xnor2_1
X_6614__108 VPWR VGND net108 sg13g2_tiehi
X_6432_ net316 VGND VPWR net864 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[10\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_2
X_3644_ _0697_ _0679_ _0696_ VPWR VGND sg13g2_nand2_1
X_3575_ _0630_ _0631_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[1\] u_angle_cordic_12b_pmod.u_vga_top.vsync
+ VPWR VGND _0632_ sg13g2_nand4_1
X_6363_ net375 _2917_ _2918_ _0513_ VPWR VGND sg13g2_nor3_1
X_5314_ _2071_ net970 net1008 VPWR VGND sg13g2_nand2_1
X_6294_ _2890_ net444 _2889_ VPWR VGND sg13g2_nand2_1
X_5245_ _2016_ _2018_ _0283_ VPWR VGND sg13g2_nor2_1
Xhold28 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[8\] VPWR VGND net785
+ sg13g2_dlygate4sd3_1
Xhold17 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[1\] VPWR VGND net774
+ sg13g2_dlygate4sd3_1
X_5176_ net380 net1408 _1959_ VPWR VGND sg13g2_xor2_1
X_6637__85 VPWR VGND net85 sg13g2_tiehi
Xhold39 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[7\] VPWR VGND net796
+ sg13g2_dlygate4sd3_1
X_4127_ _1089_ _1091_ _1094_ VPWR VGND sg13g2_nor2_1
XFILLER_28_126 VPWR VGND sg13g2_fill_2
XFILLER_43_107 VPWR VGND sg13g2_fill_2
X_4058_ _1044_ VPWR _0066_ VGND net372 _1048_ sg13g2_o21ai_1
XFILLER_45_49 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_63_clk clknet_4_2_0_clk clknet_leaf_63_clk VPWR VGND sg13g2_buf_8
XFILLER_24_343 VPWR VGND sg13g2_fill_2
XFILLER_4_748 VPWR VGND sg13g2_decap_8
XFILLER_3_258 VPWR VGND sg13g2_fill_1
XFILLER_0_976 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_54_clk clknet_4_8_0_clk clknet_leaf_54_clk VPWR VGND sg13g2_buf_8
XFILLER_30_313 VPWR VGND sg13g2_fill_2
XFILLER_30_357 VPWR VGND sg13g2_fill_1
Xhold509 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[4\] VPWR VGND net1266
+ sg13g2_dlygate4sd3_1
X_5030_ _0239_ net470 _1846_ _1847_ VPWR VGND sg13g2_and3_1
XFILLER_2_291 VPWR VGND sg13g2_fill_2
XFILLER_38_468 VPWR VGND sg13g2_fill_2
X_6634__88 VPWR VGND net88 sg13g2_tiehi
X_5932_ _2589_ net1455 _2594_ VPWR VGND sg13g2_nor2_1
XFILLER_25_129 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_45_clk clknet_4_12_0_clk clknet_leaf_45_clk VPWR VGND sg13g2_buf_8
X_5863_ _2535_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[9\]
+ _2534_ VPWR VGND sg13g2_xnor2_1
X_5794_ _2473_ net1015 _0376_ VPWR VGND sg13g2_nor2_1
XFILLER_21_324 VPWR VGND sg13g2_fill_1
XFILLER_33_195 VPWR VGND sg13g2_fill_2
X_4814_ net426 net1238 _1667_ _0203_ VPWR VGND sg13g2_nor3_1
X_4745_ VGND VPWR _1603_ _1608_ _1610_ _1607_ sg13g2_a21oi_1
X_4676_ VGND VPWR _1548_ _1550_ _1552_ _1547_ sg13g2_a21oi_1
X_6415_ net350 VGND VPWR _0024_ u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[4\] clknet_leaf_66_clk
+ sg13g2_dfrbpq_2
X_3627_ VGND VPWR _0670_ _0675_ _0680_ _0674_ sg13g2_a21oi_1
Xoutput18 net18 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_1_707 VPWR VGND sg13g2_decap_8
X_6346_ _0507_ net378 _2906_ _2907_ VPWR VGND sg13g2_and3_1
X_3558_ net919 net450 _0523_ VPWR VGND sg13g2_and2_1
X_6277_ net444 VPWR _2878_ VGND _2873_ _2877_ sg13g2_o21ai_1
X_3489_ _0559_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[7\]
+ VPWR VGND sg13g2_inv_2
XFILLER_5_1003 VPWR VGND sg13g2_decap_8
X_5228_ _2004_ net492 _2002_ VPWR VGND sg13g2_nand2_1
X_5159_ _1942_ VPWR _1945_ VGND _0569_ net380 sg13g2_o21ai_1
Xclkbuf_leaf_36_clk clknet_4_12_0_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
XFILLER_13_814 VPWR VGND sg13g2_fill_1
XFILLER_8_328 VPWR VGND sg13g2_fill_1
XFILLER_4_545 VPWR VGND sg13g2_fill_2
XFILLER_0_773 VPWR VGND sg13g2_decap_8
X_6604__118 VPWR VGND net118 sg13g2_tiehi
Xclkbuf_leaf_27_clk clknet_4_7_0_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
X_4530_ net499 VPWR _1432_ VGND _1430_ _1431_ sg13g2_o21ai_1
XFILLER_8_895 VPWR VGND sg13g2_decap_8
Xhold306 _1966_ VPWR VGND net1063 sg13g2_dlygate4sd3_1
Xhold317 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[2\] VPWR VGND net1074
+ sg13g2_dlygate4sd3_1
X_4461_ _1373_ _1362_ _1372_ VPWR VGND sg13g2_nand2_1
X_6200_ net454 VPWR _2818_ VGND _2815_ _2817_ sg13g2_o21ai_1
Xhold328 _0369_ VPWR VGND net1085 sg13g2_dlygate4sd3_1
Xhold339 _0292_ VPWR VGND net1096 sg13g2_dlygate4sd3_1
X_6131_ _2755_ _2751_ _2754_ _2757_ VPWR VGND sg13g2_a21o_1
X_4392_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[9\] _1312_ net410
+ _1314_ VPWR VGND sg13g2_nand3_1
X_6062_ _2689_ _2697_ _2698_ VPWR VGND sg13g2_and2_1
X_5013_ _1829_ VPWR _1832_ VGND _1825_ _1830_ sg13g2_o21ai_1
Xclkbuf_leaf_18_clk clknet_4_5_0_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
X_5915_ net1248 _2577_ _2579_ VPWR VGND sg13g2_nor2_1
X_6895_ net730 VGND VPWR _0523_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[2\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_1
X_5846_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[6\] net413
+ _2513_ _2520_ VPWR VGND sg13g2_a21o_1
XFILLER_21_143 VPWR VGND sg13g2_fill_1
XFILLER_22_666 VPWR VGND sg13g2_fill_2
X_5777_ net1487 net519 _2462_ VPWR VGND sg13g2_xor2_1
X_4728_ VGND VPWR _1591_ _1594_ _0189_ _1595_ sg13g2_a21oi_1
X_4659_ net432 _1536_ net1190 _0178_ VPWR VGND sg13g2_nor3_1
X_6329_ net469 net839 _0500_ VPWR VGND sg13g2_and2_1
XFILLER_29_232 VPWR VGND sg13g2_fill_2
XFILLER_26_972 VPWR VGND sg13g2_decap_8
XFILLER_16_84 VPWR VGND sg13g2_fill_1
XFILLER_9_659 VPWR VGND sg13g2_fill_2
XFILLER_5_821 VPWR VGND sg13g2_decap_8
XFILLER_5_898 VPWR VGND sg13g2_decap_8
XFILLER_4_397 VPWR VGND sg13g2_fill_2
XFILLER_17_983 VPWR VGND sg13g2_decap_8
X_3961_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[5\] VPWR _0962_
+ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[4\] _0943_ sg13g2_o21ai_1
X_5700_ net475 VPWR _2399_ VGND _2393_ _2398_ sg13g2_o21ai_1
X_6680_ net42 VGND VPWR _0289_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[1\]
+ clknet_leaf_36_clk sg13g2_dfrbpq_2
X_3892_ _0884_ _0911_ net1003 _0914_ VPWR VGND sg13g2_nand3_1
X_5631_ VGND VPWR _2334_ _2338_ _2340_ net431 sg13g2_a21oi_1
XFILLER_32_997 VPWR VGND sg13g2_fill_2
X_5562_ net515 _2278_ _2279_ VPWR VGND sg13g2_nor2_1
X_4513_ net384 net1332 _1418_ VPWR VGND sg13g2_xor2_1
XFILLER_8_681 VPWR VGND sg13g2_fill_2
Xhold103 _0635_ VPWR VGND net860 sg13g2_dlygate4sd3_1
Xhold114 _0018_ VPWR VGND net871 sg13g2_dlygate4sd3_1
X_5493_ net479 VPWR _2225_ VGND _2223_ _2224_ sg13g2_o21ai_1
Xhold125 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[0\] VPWR VGND net882 sg13g2_dlygate4sd3_1
Xhold158 _0920_ VPWR VGND net915 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_4_3_0_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
Xhold136 _0852_ VPWR VGND net893 sg13g2_dlygate4sd3_1
Xhold147 _2428_ VPWR VGND net904 sg13g2_dlygate4sd3_1
X_4444_ _1353_ _1357_ _1359_ VPWR VGND sg13g2_and2_1
Xhold169 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[4\] VPWR VGND net926
+ sg13g2_dlygate4sd3_1
X_4375_ _1299_ _1300_ _1301_ VPWR VGND sg13g2_and2_1
X_6114_ _2739_ VPWR _2742_ VGND _2735_ _2740_ sg13g2_o21ai_1
X_6045_ VGND VPWR _2676_ _2681_ _2683_ _2679_ sg13g2_a21oi_1
XFILLER_2_1028 VPWR VGND sg13g2_fill_1
X_6901__552 VPWR VGND net736 sg13g2_tiehi
XFILLER_42_739 VPWR VGND sg13g2_fill_1
X_6878_ net329 VGND VPWR _0487_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[10\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_23_964 VPWR VGND sg13g2_decap_8
X_5829_ _2505_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[5\]
+ _2504_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_802 VPWR VGND sg13g2_decap_8
Xhold670 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[1\] VPWR VGND net1427
+ sg13g2_dlygate4sd3_1
X_6453__287 VPWR VGND net287 sg13g2_tiehi
Xhold681 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[2\] VPWR VGND net1438
+ sg13g2_dlygate4sd3_1
XFILLER_2_879 VPWR VGND sg13g2_decap_8
Xhold692 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[6\] VPWR
+ VGND net1449 sg13g2_dlygate4sd3_1
XFILLER_40_1001 VPWR VGND sg13g2_fill_1
XFILLER_45_500 VPWR VGND sg13g2_fill_2
XFILLER_18_714 VPWR VGND sg13g2_fill_2
XFILLER_14_920 VPWR VGND sg13g2_decap_8
XFILLER_13_430 VPWR VGND sg13g2_fill_2
XFILLER_9_423 VPWR VGND sg13g2_fill_1
XFILLER_14_997 VPWR VGND sg13g2_decap_8
X_6432__316 VPWR VGND net316 sg13g2_tiehi
XFILLER_4_32 VPWR VGND sg13g2_fill_2
X_4160_ net495 VPWR _1121_ VGND net1104 _1120_ sg13g2_o21ai_1
X_4091_ _1069_ net821 net828 _1066_ VPWR VGND sg13g2_and3_2
XFILLER_49_894 VPWR VGND sg13g2_fill_1
X_6801_ net624 VGND VPWR _0410_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[8\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_1
X_4993_ net468 VPWR _1817_ VGND _1814_ _1816_ sg13g2_o21ai_1
X_6732_ net693 VGND VPWR _0341_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[3\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3944_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[6\] _0944_ _0945_
+ VPWR VGND sg13g2_nor2b_1
X_3875_ _0884_ _0900_ _0901_ VPWR VGND sg13g2_and2_1
XFILLER_17_1025 VPWR VGND sg13g2_decap_4
X_6663_ net59 VGND VPWR _0272_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[10\]
+ clknet_leaf_49_clk sg13g2_dfrbpq_2
X_5614_ _2323_ net1334 _2325_ VPWR VGND sg13g2_xor2_1
XFILLER_20_989 VPWR VGND sg13g2_decap_8
X_6594_ net128 VGND VPWR net1239 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[5\]
+ clknet_leaf_28_clk sg13g2_dfrbpq_1
X_5545_ net811 net525 _2266_ VPWR VGND sg13g2_xor2_1
X_5476_ net430 _2209_ _2210_ _0322_ VPWR VGND sg13g2_nor3_1
X_4427_ _1345_ _1338_ _1340_ _1344_ VPWR VGND sg13g2_and3_1
Xfanout402 _2857_ net402 VPWR VGND sg13g2_buf_2
Xfanout413 _0573_ net413 VPWR VGND sg13g2_buf_8
XFILLER_48_49 VPWR VGND sg13g2_decap_8
Xfanout435 net438 net435 VPWR VGND sg13g2_buf_8
Xfanout457 net458 net457 VPWR VGND sg13g2_buf_8
Xfanout424 net428 net424 VPWR VGND sg13g2_buf_8
Xfanout446 net447 net446 VPWR VGND sg13g2_buf_1
X_4358_ net1138 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].z_sign _1287_
+ VPWR VGND sg13g2_xor2_1
Xfanout479 net480 net479 VPWR VGND sg13g2_buf_8
X_4289_ net435 _1230_ _1231_ _0114_ VPWR VGND sg13g2_nor3_1
Xfanout468 net472 net468 VPWR VGND sg13g2_buf_8
X_6028_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[0\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[1\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[2\] _2668_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_39_371 VPWR VGND sg13g2_fill_1
XFILLER_11_912 VPWR VGND sg13g2_decap_8
XFILLER_23_794 VPWR VGND sg13g2_fill_1
XFILLER_11_989 VPWR VGND sg13g2_decap_8
XFILLER_2_610 VPWR VGND sg13g2_fill_1
XFILLER_2_676 VPWR VGND sg13g2_decap_8
XFILLER_18_588 VPWR VGND sg13g2_decap_4
XFILLER_33_536 VPWR VGND sg13g2_fill_2
X_3660_ _0712_ _0705_ _0711_ _0713_ VPWR VGND sg13g2_a21o_1
Xclkload12 clknet_4_15_0_clk clkload12/X VPWR VGND sg13g2_buf_8
X_3591_ net547 u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[4\] u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[4\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[4\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp\[11\]
+ net545 _0644_ VPWR VGND sg13g2_mux4_1
X_5330_ _2083_ _2078_ _2085_ VPWR VGND sg13g2_nor2b_1
XFILLER_6_993 VPWR VGND sg13g2_decap_8
X_5261_ _2023_ _2024_ _2028_ _2031_ VPWR VGND sg13g2_or3_1
X_4212_ _1166_ net1183 net382 VPWR VGND sg13g2_xnor2_1
X_5192_ _1971_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[5\]\[2\] _1972_
+ VPWR VGND sg13g2_nor2b_1
X_4143_ VGND VPWR _1108_ _1107_ _1106_ sg13g2_or2_1
XFILLER_28_308 VPWR VGND sg13g2_fill_1
X_4074_ _1056_ VPWR _0072_ VGND net373 _1057_ sg13g2_o21ai_1
XFILLER_49_680 VPWR VGND sg13g2_fill_2
XFILLER_36_330 VPWR VGND sg13g2_fill_1
X_6715_ net710 VGND VPWR _0324_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[6\]
+ clknet_leaf_48_clk sg13g2_dfrbpq_2
X_4976_ VGND VPWR _1800_ _1801_ _1803_ net426 sg13g2_a21oi_1
X_3927_ _0928_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[4\] _0929_
+ VPWR VGND sg13g2_nor2b_1
X_3858_ net441 VPWR _0889_ VGND net1030 _0886_ sg13g2_o21ai_1
Xclkload6 clknet_4_9_0_clk clkload6/X VPWR VGND sg13g2_buf_8
X_6646_ net76 VGND VPWR _0255_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[7\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
X_6577_ net145 VGND VPWR net1440 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[2\]
+ clknet_leaf_34_clk sg13g2_dfrbpq_1
X_3789_ VPWR VGND net914 _0835_ _0552_ _0535_ _0836_ net909 sg13g2_a221oi_1
X_5528_ _2251_ VPWR _2252_ VGND net523 _0561_ sg13g2_o21ai_1
X_6888__296 VPWR VGND net296 sg13g2_tiehi
X_5459_ _2196_ net1388 _2195_ VPWR VGND sg13g2_nand2_1
XFILLER_19_319 VPWR VGND sg13g2_fill_1
XFILLER_24_40 VPWR VGND sg13g2_fill_2
XFILLER_24_73 VPWR VGND sg13g2_fill_2
XFILLER_7_746 VPWR VGND sg13g2_decap_8
XFILLER_7_735 VPWR VGND sg13g2_fill_2
XFILLER_11_786 VPWR VGND sg13g2_fill_2
XFILLER_3_941 VPWR VGND sg13g2_decap_8
XFILLER_45_182 VPWR VGND sg13g2_fill_2
X_4830_ _1681_ net1137 net392 VPWR VGND sg13g2_xnor2_1
X_4761_ net488 VPWR _1623_ VGND _1621_ _1622_ sg13g2_o21ai_1
X_3712_ _0765_ _0763_ _0748_ VPWR VGND sg13g2_nand2b_1
X_6500_ net222 VGND VPWR net992 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[1\]
+ clknet_leaf_47_clk sg13g2_dfrbpq_1
X_4692_ _1564_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[0\]
+ net537 VPWR VGND sg13g2_nand2b_1
X_6431_ net318 VGND VPWR net1002 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[9\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_2
X_3643_ _0696_ _0667_ _0695_ VPWR VGND sg13g2_xnor2_1
X_6362_ net981 _2915_ _2918_ VPWR VGND sg13g2_nor2_1
XFILLER_6_790 VPWR VGND sg13g2_decap_8
X_3574_ _0632_ net978 net920 VPWR VGND sg13g2_nand2_1
X_5313_ VGND VPWR _0564_ net837 _0299_ _2070_ sg13g2_a21oi_1
X_6293_ _2889_ _2872_ _2887_ VPWR VGND sg13g2_nand2_1
X_5244_ _2018_ net492 _2017_ VPWR VGND sg13g2_nand2_1
X_5175_ VGND VPWR _1952_ _1955_ _1958_ _1957_ sg13g2_a21oi_1
Xhold18 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[5\] VPWR VGND net775
+ sg13g2_dlygate4sd3_1
Xhold29 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[4\] VPWR VGND net786
+ sg13g2_dlygate4sd3_1
X_4126_ net436 _1092_ _1093_ _0089_ VPWR VGND sg13g2_nor3_1
X_4057_ _1048_ _1045_ _1047_ VPWR VGND sg13g2_xnor2_1
X_4959_ _1784_ _1776_ _1788_ VPWR VGND _1780_ sg13g2_nand3b_1
X_6629_ net93 VGND VPWR net1490 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[2\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_4_727 VPWR VGND sg13g2_decap_8
XFILLER_0_955 VPWR VGND sg13g2_decap_8
XFILLER_47_403 VPWR VGND sg13g2_fill_1
XFILLER_19_105 VPWR VGND sg13g2_fill_2
XFILLER_28_661 VPWR VGND sg13g2_fill_1
XFILLER_27_182 VPWR VGND sg13g2_fill_1
XFILLER_20_1010 VPWR VGND sg13g2_decap_8
X_5931_ _2593_ net1454 _2591_ VPWR VGND sg13g2_xnor2_1
XFILLER_19_683 VPWR VGND sg13g2_fill_1
X_6620__102 VPWR VGND net102 sg13g2_tiehi
XFILLER_18_171 VPWR VGND sg13g2_fill_2
X_5862_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[8\] net413
+ _2526_ _2534_ VPWR VGND sg13g2_a21o_1
X_5793_ net457 VPWR _2474_ VGND net1014 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[0\]
+ sg13g2_o21ai_1
XFILLER_21_314 VPWR VGND sg13g2_fill_1
X_4813_ _1667_ _1661_ _1664_ _1665_ VPWR VGND sg13g2_and3_1
X_4744_ _1607_ _1608_ _1603_ _1609_ VPWR VGND sg13g2_nand3_1
XFILLER_21_347 VPWR VGND sg13g2_fill_2
X_4675_ _1551_ _1547_ _1548_ _1550_ VPWR VGND sg13g2_and3_1
X_6414_ net352 VGND VPWR net938 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[3\] clknet_leaf_66_clk
+ sg13g2_dfrbpq_1
X_3626_ _0678_ _0661_ _0677_ _0679_ VPWR VGND sg13g2_a21o_2
Xoutput19 net19 uo_out[1] VPWR VGND sg13g2_buf_1
X_6345_ _2903_ net844 net1114 _2907_ VPWR VGND sg13g2_a21o_1
X_3557_ net840 net450 _0522_ VPWR VGND sg13g2_and2_1
X_6276_ _2877_ _0543_ _2876_ VPWR VGND sg13g2_xnor2_1
X_3488_ VPWR _0558_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[6\] VGND
+ sg13g2_inv_1
X_5227_ _1993_ _2000_ _2001_ _2003_ VPWR VGND sg13g2_nor3_1
X_5158_ _1944_ net1289 _1934_ VPWR VGND sg13g2_xnor2_1
X_5089_ net478 VPWR _1884_ VGND net1033 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[0\]
+ sg13g2_o21ai_1
XFILLER_29_447 VPWR VGND sg13g2_fill_1
X_4109_ VGND VPWR _1080_ _1079_ _1077_ sg13g2_or2_1
XFILLER_25_675 VPWR VGND sg13g2_fill_2
XFILLER_0_752 VPWR VGND sg13g2_decap_8
XFILLER_8_874 VPWR VGND sg13g2_decap_8
XFILLER_7_351 VPWR VGND sg13g2_fill_1
Xhold307 _0276_ VPWR VGND net1064 sg13g2_dlygate4sd3_1
X_4460_ net387 VPWR _1372_ VGND net1158 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[4\]
+ sg13g2_o21ai_1
Xhold318 _0328_ VPWR VGND net1075 sg13g2_dlygate4sd3_1
Xhold329 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[8\] VPWR VGND net1086
+ sg13g2_dlygate4sd3_1
X_4391_ _1312_ net410 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[9\]
+ _1313_ VPWR VGND sg13g2_a21o_1
X_6130_ VGND VPWR _2751_ _2755_ _0430_ _2756_ sg13g2_a21oi_1
X_6061_ _2697_ net416 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[6\]
+ VPWR VGND sg13g2_nand2_1
X_5012_ VGND VPWR _1825_ _1830_ _0237_ _1831_ sg13g2_a21oi_1
XFILLER_38_266 VPWR VGND sg13g2_fill_2
X_5914_ _2578_ net1248 _2577_ VPWR VGND sg13g2_nand2_1
X_6894_ net729 VGND VPWR _0522_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[1\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_35_984 VPWR VGND sg13g2_fill_1
X_5845_ VGND VPWR _2512_ _2517_ _2519_ _2515_ sg13g2_a21oi_1
X_6630__92 VPWR VGND net92 sg13g2_tiehi
XFILLER_35_995 VPWR VGND sg13g2_fill_2
X_5776_ net519 net1487 _2461_ VPWR VGND sg13g2_nor2b_1
X_4727_ net488 VPWR _1595_ VGND _1591_ _1594_ sg13g2_o21ai_1
X_4658_ VGND VPWR _1531_ _1533_ _1537_ _1535_ sg13g2_a21oi_1
X_3609_ VGND VPWR net409 net408 _0662_ net407 sg13g2_a21oi_1
X_4589_ VPWR VGND _1477_ _1478_ _1467_ _0608_ _1479_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[7\]
+ sg13g2_a221oi_1
XFILLER_27_1016 VPWR VGND sg13g2_decap_8
XFILLER_27_1027 VPWR VGND sg13g2_fill_2
X_6328_ net463 net789 _0499_ VPWR VGND sg13g2_and2_1
X_6259_ _2862_ net506 net555 VPWR VGND sg13g2_nand2_2
XFILLER_17_439 VPWR VGND sg13g2_fill_1
XFILLER_16_74 VPWR VGND sg13g2_fill_1
XFILLER_40_475 VPWR VGND sg13g2_fill_2
XFILLER_5_800 VPWR VGND sg13g2_decap_8
XFILLER_10_1020 VPWR VGND sg13g2_decap_8
X_6610__112 VPWR VGND net112 sg13g2_tiehi
XFILLER_5_877 VPWR VGND sg13g2_decap_8
XFILLER_17_962 VPWR VGND sg13g2_decap_8
X_3960_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[3\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[2\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[4\] _0960_ _0961_ VPWR VGND
+ sg13g2_nor4_1
XFILLER_35_269 VPWR VGND sg13g2_fill_2
X_3891_ VGND VPWR _0884_ _0911_ _0913_ net1003 sg13g2_a21oi_1
X_5630_ _2334_ _2338_ _2339_ VPWR VGND sg13g2_nor2_1
X_5561_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[0\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[1\]
+ _2278_ VPWR VGND sg13g2_nor2_1
X_4512_ net1332 net384 _1417_ VPWR VGND sg13g2_and2_1
XFILLER_8_671 VPWR VGND sg13g2_fill_1
X_5492_ _2206_ net1285 _2224_ VPWR VGND sg13g2_xor2_1
Xhold115 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[10\] VPWR
+ VGND net872 sg13g2_dlygate4sd3_1
Xhold104 _0002_ VPWR VGND net861 sg13g2_dlygate4sd3_1
Xhold126 _0848_ VPWR VGND net883 sg13g2_dlygate4sd3_1
Xhold159 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[16\] VPWR VGND net916
+ sg13g2_dlygate4sd3_1
Xhold137 _0014_ VPWR VGND net894 sg13g2_dlygate4sd3_1
Xhold148 _0363_ VPWR VGND net905 sg13g2_dlygate4sd3_1
X_4443_ _1358_ net1369 net386 VPWR VGND sg13g2_xnor2_1
X_4374_ net410 VPWR _1300_ VGND net1110 net1121 sg13g2_o21ai_1
X_6113_ VGND VPWR _2735_ _2740_ _0428_ _2741_ sg13g2_a21oi_1
X_6044_ VGND VPWR _2675_ net1296 _0418_ _2682_ sg13g2_a21oi_1
XFILLER_26_258 VPWR VGND sg13g2_fill_1
XFILLER_23_943 VPWR VGND sg13g2_decap_8
X_6877_ net331 VGND VPWR _0486_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[9\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_2
X_5828_ net514 _2497_ _2504_ VPWR VGND sg13g2_nor2_1
X_5759_ _2447_ net518 net1084 VPWR VGND sg13g2_nand2b_1
Xhold660 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[5\] VPWR VGND net1417
+ sg13g2_dlygate4sd3_1
XFILLER_2_858 VPWR VGND sg13g2_decap_8
Xhold671 _2477_ VPWR VGND net1428 sg13g2_dlygate4sd3_1
Xhold682 _1574_ VPWR VGND net1439 sg13g2_dlygate4sd3_1
Xhold693 _2413_ VPWR VGND net1450 sg13g2_dlygate4sd3_1
XFILLER_45_578 VPWR VGND sg13g2_fill_1
XFILLER_32_228 VPWR VGND sg13g2_fill_1
XFILLER_14_976 VPWR VGND sg13g2_decap_8
XFILLER_13_475 VPWR VGND sg13g2_fill_1
XFILLER_4_184 VPWR VGND sg13g2_fill_1
X_4090_ VGND VPWR net828 _1066_ _1068_ net821 sg13g2_a21oi_1
XFILLER_48_394 VPWR VGND sg13g2_fill_1
X_6800_ net625 VGND VPWR _0409_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[7\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_1
X_4992_ net398 net1186 _1816_ VPWR VGND sg13g2_xor2_1
X_6731_ net694 VGND VPWR net1303 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[2\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_1
XFILLER_17_1004 VPWR VGND sg13g2_decap_8
X_3943_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[4\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[5\]
+ _0943_ _0944_ VPWR VGND sg13g2_nor3_1
X_3874_ _0897_ _0898_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[9\] _0900_ VPWR VGND
+ _0899_ sg13g2_nand4_1
X_6662_ net60 VGND VPWR net1290 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[9\]
+ clknet_leaf_51_clk sg13g2_dfrbpq_2
X_5613_ net1334 _2323_ _2324_ VPWR VGND sg13g2_and2_1
XFILLER_20_968 VPWR VGND sg13g2_decap_8
X_6853__382 VPWR VGND net566 sg13g2_tiehi
X_6593_ net129 VGND VPWR _0202_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[4\]
+ clknet_leaf_26_clk sg13g2_dfrbpq_2
X_5544_ VPWR VGND _2263_ _2262_ _2260_ _0553_ _2265_ net1124 sg13g2_a221oi_1
X_5475_ _2210_ _2202_ _2205_ _2208_ VPWR VGND sg13g2_and3_1
X_4426_ _1344_ net1471 net387 VPWR VGND sg13g2_xnor2_1
Xfanout414 _0573_ net414 VPWR VGND sg13g2_buf_1
Xfanout403 _0647_ net403 VPWR VGND sg13g2_buf_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
Xfanout447 net451 net447 VPWR VGND sg13g2_buf_2
Xfanout425 net428 net425 VPWR VGND sg13g2_buf_8
X_4357_ VGND VPWR _1282_ _1284_ _0127_ _1286_ sg13g2_a21oi_1
Xfanout436 net437 net436 VPWR VGND sg13g2_buf_8
Xfanout458 net461 net458 VPWR VGND sg13g2_buf_2
X_4288_ _1223_ _1229_ _1231_ VPWR VGND sg13g2_and2_1
Xfanout469 net471 net469 VPWR VGND sg13g2_buf_8
XFILLER_46_309 VPWR VGND sg13g2_fill_2
X_6027_ VGND VPWR _2659_ _2663_ _2667_ _2662_ sg13g2_a21oi_1
XFILLER_42_537 VPWR VGND sg13g2_fill_1
X_6600__122 VPWR VGND net122 sg13g2_tiehi
XFILLER_11_968 VPWR VGND sg13g2_decap_8
XFILLER_7_939 VPWR VGND sg13g2_decap_8
Xhold490 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].z_sign VPWR VGND
+ net1247 sg13g2_dlygate4sd3_1
XFILLER_46_810 VPWR VGND sg13g2_fill_2
X_6700__555 VPWR VGND net739 sg13g2_tiehi
XFILLER_13_272 VPWR VGND sg13g2_fill_2
Xclkload13 clknet_leaf_66_clk clkload13/X VPWR VGND sg13g2_buf_8
X_3590_ net546 u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[5\] u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[5\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[5\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp\[11\]
+ net544 _0643_ VPWR VGND sg13g2_mux4_1
XFILLER_6_972 VPWR VGND sg13g2_decap_8
X_5260_ net430 _2029_ net1228 _0286_ VPWR VGND sg13g2_nor3_1
X_4211_ VPWR VGND net1208 _1164_ net382 net991 _1165_ _1154_ sg13g2_a221oi_1
X_6649__73 VPWR VGND net73 sg13g2_tiehi
X_5191_ _1971_ _0568_ _1970_ VPWR VGND sg13g2_xnor2_1
X_4142_ net1115 net533 _1107_ VPWR VGND sg13g2_xor2_1
X_4073_ net919 net840 net879 _1057_ VPWR VGND sg13g2_or3_1
X_6920__258 VPWR VGND net258 sg13g2_tiehi
X_4975_ _1800_ _1801_ _1802_ VPWR VGND sg13g2_nor2_1
X_6714_ net711 VGND VPWR _0323_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[5\]
+ clknet_leaf_48_clk sg13g2_dfrbpq_2
X_3926_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[3\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[2\]
+ _0927_ _0928_ VPWR VGND sg13g2_nor3_1
X_3857_ net1030 _0886_ _0888_ VPWR VGND sg13g2_and2_1
Xclkload7 clknet_4_10_0_clk clkload7/X VPWR VGND sg13g2_buf_8
X_6645_ net77 VGND VPWR _0254_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[6\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3788_ net906 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[1\] _0835_ VPWR VGND sg13g2_xor2_1
X_6576_ net146 VGND VPWR net1018 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[1\]
+ clknet_leaf_33_clk sg13g2_dfrbpq_1
XFILLER_4_909 VPWR VGND sg13g2_decap_8
X_5527_ _0332_ net481 _2250_ _2251_ VPWR VGND sg13g2_and3_1
X_5458_ _2195_ net1386 _2194_ VPWR VGND sg13g2_xnor2_1
X_5389_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[10\] _2132_ _2136_
+ VPWR VGND sg13g2_and2_1
X_4409_ _1329_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[11\] _1327_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_27_364 VPWR VGND sg13g2_fill_1
XFILLER_24_63 VPWR VGND sg13g2_fill_1
XFILLER_7_725 VPWR VGND sg13g2_fill_2
XFILLER_10_297 VPWR VGND sg13g2_fill_2
XFILLER_40_51 VPWR VGND sg13g2_fill_2
XFILLER_3_920 VPWR VGND sg13g2_decap_8
XFILLER_3_997 VPWR VGND sg13g2_decap_8
XFILLER_49_82 VPWR VGND sg13g2_decap_8
X_6646__76 VPWR VGND net76 sg13g2_tiehi
XFILLER_38_618 VPWR VGND sg13g2_fill_1
XFILLER_18_397 VPWR VGND sg13g2_fill_2
X_4760_ net400 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[11\] _1622_
+ VPWR VGND sg13g2_xor2_1
XFILLER_33_389 VPWR VGND sg13g2_fill_1
XFILLER_14_1018 VPWR VGND sg13g2_decap_8
X_3711_ _0763_ _0748_ _0764_ VPWR VGND sg13g2_nor2b_1
X_4691_ net994 _1562_ _0184_ VPWR VGND sg13g2_nor2b_1
X_6430_ net320 VGND VPWR _0039_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[8\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_2
X_3642_ _0695_ _0680_ _0693_ VPWR VGND sg13g2_xnor2_1
X_6361_ net981 _2915_ _2917_ VPWR VGND sg13g2_and2_1
X_3573_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[10\] u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[9\]
+ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[4\] _0535_ _0631_ VPWR VGND sg13g2_nor4_1
X_5312_ VGND VPWR _2068_ _2069_ _0298_ _2070_ sg13g2_a21oi_1
X_6292_ _2872_ _2887_ _2888_ VPWR VGND sg13g2_nor2_1
X_5243_ _2015_ VPWR _2017_ VGND _2010_ _2013_ sg13g2_o21ai_1
Xhold19 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[7\] VPWR VGND net776
+ sg13g2_dlygate4sd3_1
X_5174_ _1957_ _1949_ _1956_ VPWR VGND sg13g2_nand2_1
X_4125_ _1093_ _1087_ _1089_ _1091_ VPWR VGND sg13g2_and3_1
X_4056_ _1047_ net982 net548 VPWR VGND sg13g2_xnor2_1
XFILLER_43_109 VPWR VGND sg13g2_fill_1
XFILLER_24_345 VPWR VGND sg13g2_fill_1
XFILLER_36_172 VPWR VGND sg13g2_fill_1
X_4958_ _0227_ net464 net1465 _1787_ VPWR VGND sg13g2_and3_1
X_4889_ VGND VPWR _1726_ _1728_ _0216_ _1729_ sg13g2_a21oi_1
X_3909_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[9\] _0922_ _0925_ VPWR VGND sg13g2_and2_1
XFILLER_20_551 VPWR VGND sg13g2_fill_2
X_6628_ net94 VGND VPWR net1053 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[1\]
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_4_706 VPWR VGND sg13g2_decap_8
X_6559_ net163 VGND VPWR _0168_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[9\]
+ clknet_leaf_39_clk sg13g2_dfrbpq_1
XFILLER_0_934 VPWR VGND sg13g2_decap_8
XFILLER_43_610 VPWR VGND sg13g2_fill_1
X_6643__79 VPWR VGND net79 sg13g2_tiehi
XFILLER_35_51 VPWR VGND sg13g2_fill_2
XFILLER_24_890 VPWR VGND sg13g2_fill_2
XFILLER_3_794 VPWR VGND sg13g2_decap_8
X_5930_ _2591_ net1454 _2592_ VPWR VGND sg13g2_nor2b_1
XFILLER_25_109 VPWR VGND sg13g2_fill_1
X_5861_ _2529_ _2525_ _2528_ _2533_ VPWR VGND sg13g2_a21o_1
XFILLER_22_827 VPWR VGND sg13g2_fill_1
X_5792_ net1014 net1242 _2473_ VPWR VGND sg13g2_and2_1
X_4812_ VGND VPWR _1661_ _1664_ _1666_ _1665_ sg13g2_a21oi_1
X_6919__260 VPWR VGND net260 sg13g2_tiehi
X_4743_ _1604_ VPWR _1608_ VGND _1596_ _1600_ sg13g2_o21ai_1
X_6413_ net354 VGND VPWR _0022_ u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[2\] clknet_leaf_66_clk
+ sg13g2_dfrbpq_1
X_4674_ _1550_ net394 _1549_ VPWR VGND sg13g2_nand2b_1
X_3625_ _0678_ _0666_ _0676_ VPWR VGND sg13g2_xnor2_1
X_6344_ net1114 _2903_ net844 _2906_ VPWR VGND sg13g2_nand3_1
X_3556_ net879 net451 _0519_ VPWR VGND sg13g2_and2_1
X_6275_ net555 net506 _2875_ _2876_ VPWR VGND sg13g2_a21o_1
X_5226_ _2000_ VPWR _2002_ VGND _1993_ _2001_ sg13g2_o21ai_1
X_3487_ _0557_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[5\]
+ VPWR VGND sg13g2_inv_2
X_5157_ _1943_ _1942_ _0270_ VPWR VGND sg13g2_nor2b_1
X_5088_ _1883_ net1033 net1101 VPWR VGND sg13g2_nand2_1
X_4108_ _1079_ net532 net1057 VPWR VGND sg13g2_xnor2_1
X_4039_ _1032_ net548 net918 VPWR VGND sg13g2_nand2b_1
XFILLER_25_621 VPWR VGND sg13g2_fill_2
XFILLER_25_654 VPWR VGND sg13g2_fill_1
XFILLER_12_315 VPWR VGND sg13g2_fill_1
XFILLER_4_547 VPWR VGND sg13g2_fill_1
XFILLER_0_731 VPWR VGND sg13g2_decap_8
XFILLER_48_768 VPWR VGND sg13g2_fill_2
XFILLER_30_112 VPWR VGND sg13g2_fill_2
XFILLER_8_853 VPWR VGND sg13g2_decap_8
XFILLER_12_893 VPWR VGND sg13g2_decap_8
Xhold308 net22 VPWR VGND net1065 sg13g2_dlygate4sd3_1
Xhold319 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[0\] VPWR
+ VGND net1076 sg13g2_dlygate4sd3_1
X_4390_ VGND VPWR _1312_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[8\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[7\] sg13g2_or2_1
XFILLER_3_591 VPWR VGND sg13g2_fill_1
X_6060_ net1523 _2696_ _0420_ VPWR VGND sg13g2_and2_1
X_5011_ net469 VPWR _1831_ VGND _1825_ _1830_ sg13g2_o21ai_1
X_5913_ _2577_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[6\] _2576_
+ VPWR VGND sg13g2_xnor2_1
X_6893_ net728 VGND VPWR _0519_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[0\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_1
X_5844_ VGND VPWR _2511_ net1307 _0382_ _2518_ sg13g2_a21oi_1
XFILLER_22_668 VPWR VGND sg13g2_fill_1
XFILLER_21_178 VPWR VGND sg13g2_fill_1
XFILLER_22_679 VPWR VGND sg13g2_fill_1
X_5775_ _2456_ _2458_ _2460_ VPWR VGND sg13g2_and2_1
X_4726_ net401 net1293 _1594_ VPWR VGND sg13g2_xor2_1
X_4657_ _1536_ _1531_ _1533_ _1535_ VPWR VGND sg13g2_and3_1
Xhold820 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[0\] VPWR VGND net1577 sg13g2_dlygate4sd3_1
X_3608_ _0661_ net409 net408 net407 VPWR VGND sg13g2_and3_2
X_4588_ _1478_ _1470_ _1468_ VPWR VGND sg13g2_nand2b_1
X_6327_ net462 net794 _0498_ VPWR VGND sg13g2_and2_1
X_3539_ VPWR _0609_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[2\]
+ VGND sg13g2_inv_1
X_6258_ VGND VPWR _2860_ _2861_ _0453_ net421 sg13g2_a21oi_1
X_5209_ _1985_ net1380 _1987_ VPWR VGND sg13g2_xor2_1
X_6189_ _2804_ _2800_ _2803_ _2808_ VPWR VGND sg13g2_a21o_1
XFILLER_18_919 VPWR VGND sg13g2_decap_8
XFILLER_29_256 VPWR VGND sg13g2_fill_1
XFILLER_38_790 VPWR VGND sg13g2_fill_1
XFILLER_41_922 VPWR VGND sg13g2_fill_2
XFILLER_5_856 VPWR VGND sg13g2_decap_8
XFILLER_17_941 VPWR VGND sg13g2_decap_8
X_3890_ _0885_ net978 _0912_ _0034_ VPWR VGND sg13g2_a21o_1
XFILLER_31_421 VPWR VGND sg13g2_fill_2
X_5560_ VGND VPWR _2268_ _2273_ _2277_ _2272_ sg13g2_a21oi_1
XFILLER_31_498 VPWR VGND sg13g2_decap_8
X_5491_ _2214_ _2221_ _2222_ _2223_ VPWR VGND sg13g2_nor3_1
X_4511_ _1410_ net543 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[10\]
+ _1416_ VPWR VGND sg13g2_mux2_1
Xhold116 _0183_ VPWR VGND net873 sg13g2_dlygate4sd3_1
Xhold105 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[3\] VPWR VGND net862
+ sg13g2_dlygate4sd3_1
X_4442_ _0141_ net486 _1356_ _1357_ VPWR VGND sg13g2_and3_1
Xhold138 net21 VPWR VGND net895 sg13g2_dlygate4sd3_1
Xhold149 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[1\] VPWR VGND net906 sg13g2_dlygate4sd3_1
Xhold127 _0012_ VPWR VGND net884 sg13g2_dlygate4sd3_1
X_4373_ _1299_ _1297_ _1294_ VPWR VGND sg13g2_nand2b_1
X_6112_ net452 VPWR _2741_ VGND _2735_ _2740_ sg13g2_o21ai_1
X_6043_ net452 VPWR _2682_ VGND _2675_ _2680_ sg13g2_o21ai_1
XFILLER_2_1019 VPWR VGND sg13g2_decap_8
XFILLER_23_922 VPWR VGND sg13g2_decap_8
X_6876_ net333 VGND VPWR _0485_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[8\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_1
X_5827_ _2500_ VPWR _2503_ VGND _2495_ _2501_ sg13g2_o21ai_1
XFILLER_23_999 VPWR VGND sg13g2_decap_8
X_5758_ _2442_ VPWR _2446_ VGND _2443_ _2444_ sg13g2_o21ai_1
X_4709_ _1579_ net1311 _1578_ VPWR VGND sg13g2_nand2b_1
X_5689_ net1456 _2388_ _2389_ VPWR VGND sg13g2_and2_1
Xhold650 _0432_ VPWR VGND net1407 sg13g2_dlygate4sd3_1
Xhold672 _0378_ VPWR VGND net1429 sg13g2_dlygate4sd3_1
XFILLER_2_837 VPWR VGND sg13g2_decap_8
Xhold661 _0305_ VPWR VGND net1418 sg13g2_dlygate4sd3_1
Xhold683 _0186_ VPWR VGND net1440 sg13g2_dlygate4sd3_1
XFILLER_1_358 VPWR VGND sg13g2_fill_1
Xhold694 _0360_ VPWR VGND net1451 sg13g2_dlygate4sd3_1
XFILLER_26_760 VPWR VGND sg13g2_fill_2
XFILLER_13_432 VPWR VGND sg13g2_fill_1
XFILLER_14_955 VPWR VGND sg13g2_decap_8
XFILLER_48_351 VPWR VGND sg13g2_fill_1
X_4991_ _1815_ net1186 net398 VPWR VGND sg13g2_nand2_1
X_6730_ net695 VGND VPWR net1232 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[1\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3942_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt_sum\[5\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[1\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[2\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[3\]
+ _0943_ VPWR VGND sg13g2_or4_1
X_3873_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[4\] u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[1\]
+ _0632_ _0899_ VPWR VGND sg13g2_nor3_1
X_6661_ net61 VGND VPWR _0270_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[8\]
+ clknet_leaf_49_clk sg13g2_dfrbpq_2
X_6592_ net130 VGND VPWR _0201_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[3\]
+ clknet_leaf_26_clk sg13g2_dfrbpq_2
X_5612_ _2323_ _0597_ _2322_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_947 VPWR VGND sg13g2_decap_8
XFILLER_32_796 VPWR VGND sg13g2_fill_2
XFILLER_9_981 VPWR VGND sg13g2_decap_8
X_5543_ VGND VPWR _2261_ net1172 _0335_ _2264_ sg13g2_a21oi_1
X_5474_ VGND VPWR _2202_ _2205_ _2209_ _2208_ sg13g2_a21oi_1
X_4425_ net1471 net387 _1343_ VPWR VGND sg13g2_and2_1
X_4356_ _1286_ net503 _1285_ VPWR VGND sg13g2_nand2_1
Xfanout404 _0646_ net404 VPWR VGND sg13g2_buf_8
XFILLER_24_1009 VPWR VGND sg13g2_decap_8
Xfanout426 net428 net426 VPWR VGND sg13g2_buf_8
Xfanout415 _0564_ net415 VPWR VGND sg13g2_buf_8
Xfanout448 net449 net448 VPWR VGND sg13g2_buf_2
Xfanout437 net438 net437 VPWR VGND sg13g2_buf_8
Xfanout459 net461 net459 VPWR VGND sg13g2_buf_8
X_4287_ _1223_ _1229_ _1230_ VPWR VGND sg13g2_nor2_1
X_6860__365 VPWR VGND net365 sg13g2_tiehi
X_6026_ _2665_ _2666_ _0416_ VPWR VGND sg13g2_nor2b_1
X_6859_ net367 VGND VPWR _0468_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[3\]
+ clknet_leaf_64_clk sg13g2_dfrbpq_1
XFILLER_23_763 VPWR VGND sg13g2_fill_2
XFILLER_11_947 VPWR VGND sg13g2_decap_8
XFILLER_22_262 VPWR VGND sg13g2_fill_2
XFILLER_7_918 VPWR VGND sg13g2_decap_8
Xheichips25_CORDIC_573 VPWR VGND uio_oe[7] sg13g2_tiehi
XFILLER_13_98 VPWR VGND sg13g2_fill_2
Xhold480 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[4\] VPWR VGND net1237
+ sg13g2_dlygate4sd3_1
Xhold491 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[2\] VPWR
+ VGND net1248 sg13g2_dlygate4sd3_1
XFILLER_46_855 VPWR VGND sg13g2_fill_2
X_6499__223 VPWR VGND net223 sg13g2_tiehi
XFILLER_6_951 VPWR VGND sg13g2_decap_8
X_4210_ _1151_ _1156_ _1160_ _1164_ VPWR VGND sg13g2_nor3_1
X_5190_ net527 _1969_ _1970_ VPWR VGND sg13g2_nor2_1
X_4141_ _1095_ _1104_ _1105_ _1106_ VPWR VGND sg13g2_nor3_1
XFILLER_49_660 VPWR VGND sg13g2_fill_2
XFILLER_23_1020 VPWR VGND sg13g2_decap_8
X_4072_ _1056_ _0523_ _1054_ VPWR VGND sg13g2_nand2_1
X_6408__364 VPWR VGND net364 sg13g2_tiehi
X_4974_ _1801_ net1122 net397 VPWR VGND sg13g2_xnor2_1
X_3925_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[1\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[0\]
+ _0927_ VPWR VGND sg13g2_and2_1
X_6713_ net712 VGND VPWR net1503 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[4\]
+ clknet_leaf_48_clk sg13g2_dfrbpq_2
X_6644_ net78 VGND VPWR _0253_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[5\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
Xclkload8 clknet_4_11_0_clk clkload8/X VPWR VGND sg13g2_buf_8
X_3856_ _0886_ _0887_ _0025_ VPWR VGND sg13g2_nor2_1
X_3787_ net869 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[7\] _0834_ VPWR VGND sg13g2_xor2_1
XFILLER_30_1013 VPWR VGND sg13g2_decap_8
X_6575_ net147 VGND VPWR net995 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[0\]
+ clknet_leaf_33_clk sg13g2_dfrbpq_1
X_5526_ _2248_ VPWR _2251_ VGND _2245_ _2249_ sg13g2_o21ai_1
X_5457_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[10\] net418 _2187_
+ _2194_ VPWR VGND sg13g2_a21o_1
X_4408_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[11\] _1327_ _1328_
+ VPWR VGND sg13g2_nor2_1
XFILLER_8_1014 VPWR VGND sg13g2_decap_8
X_5388_ VGND VPWR _2131_ _2134_ _0309_ _2135_ sg13g2_a21oi_1
X_4339_ _0124_ net502 _1270_ _1271_ VPWR VGND sg13g2_and3_1
X_6009_ _2652_ net1046 net1076 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_66_clk clknet_4_0_0_clk clknet_leaf_66_clk VPWR VGND sg13g2_buf_8
XFILLER_24_42 VPWR VGND sg13g2_fill_1
XFILLER_7_737 VPWR VGND sg13g2_fill_1
XFILLER_6_247 VPWR VGND sg13g2_fill_1
XFILLER_6_0 VPWR VGND sg13g2_fill_1
XFILLER_3_976 VPWR VGND sg13g2_decap_8
XFILLER_2_464 VPWR VGND sg13g2_fill_2
XFILLER_49_61 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_57_clk clknet_4_8_0_clk clknet_leaf_57_clk VPWR VGND sg13g2_buf_8
XFILLER_45_184 VPWR VGND sg13g2_fill_1
XFILLER_14_582 VPWR VGND sg13g2_decap_4
X_3710_ _0763_ _0681_ _0761_ VPWR VGND sg13g2_xnor2_1
X_4690_ net482 VPWR _1563_ VGND net993 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[0\]
+ sg13g2_o21ai_1
X_3641_ _0680_ _0693_ _0694_ VPWR VGND sg13g2_nor2b_1
X_3572_ net914 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[7\] u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[6\]
+ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[5\] _0630_ VPWR VGND sg13g2_and4_1
X_6360_ net375 _2915_ _2916_ _0512_ VPWR VGND sg13g2_nor3_1
X_5311_ net496 VPWR _2070_ VGND _2068_ _2069_ sg13g2_o21ai_1
X_6291_ _2887_ _2882_ _2885_ VPWR VGND sg13g2_nand2_1
X_5242_ _2010_ _2013_ _2015_ _2016_ VPWR VGND sg13g2_nor3_1
X_5173_ _1935_ VPWR _1956_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[10\]
+ net1291 sg13g2_o21ai_1
XFILLER_39_0 VPWR VGND sg13g2_fill_2
X_4124_ VGND VPWR _1087_ _1089_ _1092_ _1091_ sg13g2_a21oi_1
Xinput1 rst_n net1 VPWR VGND sg13g2_buf_2
Xclkbuf_leaf_48_clk clknet_4_11_0_clk clknet_leaf_48_clk VPWR VGND sg13g2_buf_8
X_4055_ VGND VPWR _1046_ net548 net982 sg13g2_or2_1
X_4957_ _1782_ _1779_ _1785_ _1787_ VPWR VGND sg13g2_a21o_1
X_4888_ net485 VPWR _1729_ VGND _1726_ _1728_ sg13g2_o21ai_1
X_3908_ _0923_ VPWR _0040_ VGND _0909_ _0924_ sg13g2_o21ai_1
X_3839_ VGND VPWR net554 net857 _0875_ net874 sg13g2_a21oi_1
X_6627_ net95 VGND VPWR net990 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[0\]
+ clknet_leaf_27_clk sg13g2_dfrbpq_1
X_6558_ net164 VGND VPWR net1088 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[8\]
+ clknet_leaf_39_clk sg13g2_dfrbpq_1
X_6489_ net233 VGND VPWR _0098_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[3\]
+ clknet_leaf_50_clk sg13g2_dfrbpq_2
X_5509_ VPWR _2237_ _2236_ VGND sg13g2_inv_1
XFILLER_0_913 VPWR VGND sg13g2_decap_8
X_6489__233 VPWR VGND net233 sg13g2_tiehi
XFILLER_19_107 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_39_clk clknet_4_15_0_clk clknet_leaf_39_clk VPWR VGND sg13g2_buf_8
XFILLER_16_803 VPWR VGND sg13g2_fill_1
XFILLER_27_162 VPWR VGND sg13g2_fill_2
XFILLER_42_110 VPWR VGND sg13g2_fill_2
XFILLER_27_173 VPWR VGND sg13g2_fill_1
X_6496__226 VPWR VGND net226 sg13g2_tiehi
XFILLER_11_563 VPWR VGND sg13g2_fill_2
XFILLER_3_773 VPWR VGND sg13g2_decap_8
X_5860_ _0384_ net458 _2531_ _2532_ VPWR VGND sg13g2_and3_1
X_6642__80 VPWR VGND net80 sg13g2_tiehi
X_4811_ _1665_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[5\] net391
+ VPWR VGND sg13g2_xnor2_1
X_5791_ VGND VPWR _0592_ net826 _0375_ _2472_ sg13g2_a21oi_1
X_4742_ _1607_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[8\] _1592_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_21_349 VPWR VGND sg13g2_fill_1
X_4673_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[0\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[1\]
+ _1549_ VPWR VGND sg13g2_nor2_1
X_6412_ net356 VGND VPWR net876 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[1\] clknet_leaf_66_clk
+ sg13g2_dfrbpq_1
X_3624_ _0666_ _0676_ _0677_ VPWR VGND sg13g2_nor2b_1
X_3555_ VPWR _0625_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[10\]
+ VGND sg13g2_inv_1
X_6343_ VGND VPWR net844 _2903_ _0506_ _2905_ sg13g2_a21oi_1
X_3486_ VPWR _0556_ net1517 VGND sg13g2_inv_1
X_6274_ net506 net555 _2874_ _2875_ VPWR VGND sg13g2_nor3_1
X_5225_ VPWR VGND net1542 _1986_ _1992_ _1983_ _2001_ _1987_ sg13g2_a221oi_1
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_1017 VPWR VGND sg13g2_decap_8
X_5156_ net493 VPWR _1943_ VGND _1940_ _1941_ sg13g2_o21ai_1
X_4107_ _1078_ net532 net1057 VPWR VGND sg13g2_nand2_1
X_5087_ net803 net423 _0261_ VPWR VGND sg13g2_nor2_1
XFILLER_44_419 VPWR VGND sg13g2_fill_2
XFILLER_38_972 VPWR VGND sg13g2_fill_2
X_4038_ _1031_ net918 net376 VPWR VGND sg13g2_nand2_1
XFILLER_25_677 VPWR VGND sg13g2_fill_1
XFILLER_24_165 VPWR VGND sg13g2_fill_1
X_5989_ VGND VPWR _2637_ _2636_ _2634_ sg13g2_or2_1
XFILLER_21_76 VPWR VGND sg13g2_fill_2
XFILLER_0_710 VPWR VGND sg13g2_decap_8
XFILLER_43_1001 VPWR VGND sg13g2_fill_1
XFILLER_0_787 VPWR VGND sg13g2_decap_8
X_6463__269 VPWR VGND net269 sg13g2_tiehi
XFILLER_8_832 VPWR VGND sg13g2_decap_8
XFILLER_12_872 VPWR VGND sg13g2_decap_8
Xhold309 _0830_ VPWR VGND net1066 sg13g2_dlygate4sd3_1
XFILLER_30_4 VPWR VGND sg13g2_fill_1
X_5010_ _1830_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[1\] _1828_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_26_419 VPWR VGND sg13g2_fill_2
XFILLER_38_268 VPWR VGND sg13g2_fill_1
XFILLER_47_780 VPWR VGND sg13g2_fill_1
X_5912_ net512 _2575_ _2576_ VPWR VGND sg13g2_nor2_1
X_6892_ net727 VGND VPWR net442 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.x_start\[0\]
+ clknet_leaf_0_clk sg13g2_dfrbpq_1
X_5843_ net457 VPWR _2518_ VGND _2511_ _2516_ sg13g2_o21ai_1
XFILLER_34_474 VPWR VGND sg13g2_fill_1
X_6479__243 VPWR VGND net243 sg13g2_tiehi
X_5774_ VGND VPWR _2455_ _2457_ _0371_ _2459_ sg13g2_a21oi_1
X_4725_ net1293 net401 _1593_ VPWR VGND sg13g2_nor2_1
X_4656_ _1535_ net1189 net393 VPWR VGND sg13g2_xnor2_1
Xhold810 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[7\] VPWR VGND net1567
+ sg13g2_dlygate4sd3_1
X_3607_ net409 net407 _0660_ VPWR VGND sg13g2_and2_1
X_4587_ _1471_ _1474_ _1477_ VPWR VGND sg13g2_nor2_1
X_3538_ _0608_ net540 VPWR VGND sg13g2_inv_2
X_6326_ net462 net785 _0497_ VPWR VGND sg13g2_and2_1
X_6257_ net402 _2859_ net555 _2861_ VPWR VGND sg13g2_nand3_1
X_3469_ _0539_ net554 VPWR VGND sg13g2_inv_2
X_6486__236 VPWR VGND net236 sg13g2_tiehi
X_5208_ net1380 _1985_ _1986_ VPWR VGND sg13g2_and2_1
X_6188_ VGND VPWR _2800_ _2804_ _2807_ _2803_ sg13g2_a21oi_1
X_5139_ VGND VPWR _1928_ _1927_ _1919_ sg13g2_or2_1
XFILLER_16_32 VPWR VGND sg13g2_fill_1
XFILLER_26_986 VPWR VGND sg13g2_decap_8
XFILLER_40_433 VPWR VGND sg13g2_fill_2
X_6870__345 VPWR VGND net345 sg13g2_tiehi
X_6493__229 VPWR VGND net229 sg13g2_tiehi
XFILLER_5_835 VPWR VGND sg13g2_decap_8
XFILLER_0_551 VPWR VGND sg13g2_fill_2
X_6909__282 VPWR VGND net282 sg13g2_tiehi
XFILLER_17_920 VPWR VGND sg13g2_decap_8
XFILLER_36_739 VPWR VGND sg13g2_fill_2
XFILLER_16_430 VPWR VGND sg13g2_fill_2
XFILLER_17_997 VPWR VGND sg13g2_decap_8
X_5490_ _2211_ VPWR _2222_ VGND _0559_ _2206_ sg13g2_o21ai_1
X_4510_ _1412_ VPWR _1415_ VGND _1409_ _1413_ sg13g2_o21ai_1
Xhold117 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[1\] VPWR VGND net874 sg13g2_dlygate4sd3_1
Xhold106 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[10\] VPWR VGND net863 sg13g2_dlygate4sd3_1
X_4441_ _1355_ _1349_ _1354_ _1357_ VPWR VGND sg13g2_a21o_1
Xhold139 _0820_ VPWR VGND net896 sg13g2_dlygate4sd3_1
Xhold128 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[7\] VPWR VGND
+ net885 sg13g2_dlygate4sd3_1
X_6111_ _2740_ net1076 net1265 VPWR VGND sg13g2_xnor2_1
X_4372_ VGND VPWR _1296_ _1297_ _0130_ _1298_ sg13g2_a21oi_1
X_6042_ VPWR _2681_ _2680_ VGND sg13g2_inv_1
X_6875_ net335 VGND VPWR _0484_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[7\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_34_271 VPWR VGND sg13g2_fill_2
X_5826_ VGND VPWR _2495_ _2501_ _0380_ _2502_ sg13g2_a21oi_1
XFILLER_23_978 VPWR VGND sg13g2_decap_8
X_5757_ VGND VPWR _2443_ _2444_ _0368_ _2445_ sg13g2_a21oi_1
X_4708_ _1578_ net1177 _1577_ VPWR VGND sg13g2_xnor2_1
X_6418__344 VPWR VGND net344 sg13g2_tiehi
X_5688_ _2388_ net1482 _2387_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_816 VPWR VGND sg13g2_decap_8
X_4639_ _1521_ net481 _1520_ VPWR VGND sg13g2_nand2_1
Xhold640 _0241_ VPWR VGND net1397 sg13g2_dlygate4sd3_1
Xhold662 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[3\] VPWR VGND net1419
+ sg13g2_dlygate4sd3_1
Xhold651 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[12\] VPWR VGND net1408
+ sg13g2_dlygate4sd3_1
Xhold673 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[7\] VPWR VGND net1430
+ sg13g2_dlygate4sd3_1
X_6309_ net446 net787 _0483_ VPWR VGND sg13g2_and2_1
Xhold695 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[3\] VPWR VGND net1452
+ sg13g2_dlygate4sd3_1
Xhold684 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[4\] VPWR VGND net1441
+ sg13g2_dlygate4sd3_1
XFILLER_45_525 VPWR VGND sg13g2_fill_1
XFILLER_33_709 VPWR VGND sg13g2_fill_2
XFILLER_26_772 VPWR VGND sg13g2_fill_1
XFILLER_14_934 VPWR VGND sg13g2_decap_8
XFILLER_41_720 VPWR VGND sg13g2_fill_2
XFILLER_41_764 VPWR VGND sg13g2_fill_1
XFILLER_4_153 VPWR VGND sg13g2_fill_2
XFILLER_1_882 VPWR VGND sg13g2_decap_8
XFILLER_17_750 VPWR VGND sg13g2_fill_1
X_4990_ _1811_ VPWR _1814_ VGND _1810_ _1812_ sg13g2_o21ai_1
X_3941_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt_sum\[5\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[1\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[2\] _0942_ VPWR VGND
+ sg13g2_nor3_1
X_3872_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[10\] u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[8\]
+ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[7\] _0898_ VPWR VGND sg13g2_nor3_1
X_6660_ net62 VGND VPWR _0269_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[7\]
+ clknet_leaf_50_clk sg13g2_dfrbpq_2
XFILLER_20_926 VPWR VGND sg13g2_decap_8
X_6591_ net131 VGND VPWR _0200_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[2\]
+ clknet_leaf_25_clk sg13g2_dfrbpq_2
X_5611_ net516 _2321_ _2322_ VPWR VGND sg13g2_nor2_1
X_6476__246 VPWR VGND net246 sg13g2_tiehi
XFILLER_9_960 VPWR VGND sg13g2_decap_8
X_5542_ net476 VPWR _2264_ VGND _2261_ _2263_ sg13g2_o21ai_1
XFILLER_8_481 VPWR VGND sg13g2_fill_1
X_5473_ _2208_ _0557_ _2206_ VPWR VGND sg13g2_xnor2_1
X_4424_ VGND VPWR net543 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[12\]
+ _1342_ _1335_ sg13g2_a21oi_1
Xfanout405 _0646_ net405 VPWR VGND sg13g2_buf_2
X_4355_ VGND VPWR _1285_ _1284_ _1282_ sg13g2_or2_1
Xfanout416 _0562_ net416 VPWR VGND sg13g2_buf_8
Xfanout438 net439 net438 VPWR VGND sg13g2_buf_8
Xfanout427 net428 net427 VPWR VGND sg13g2_buf_1
X_4286_ VPWR _1229_ _1228_ VGND sg13g2_inv_1
Xfanout449 net450 net449 VPWR VGND sg13g2_buf_8
X_6025_ VGND VPWR _2659_ _2664_ _2666_ net422 sg13g2_a21oi_1
XFILLER_27_503 VPWR VGND sg13g2_fill_1
XFILLER_27_514 VPWR VGND sg13g2_fill_1
X_6483__239 VPWR VGND net239 sg13g2_tiehi
XFILLER_39_385 VPWR VGND sg13g2_fill_2
X_6858_ net369 VGND VPWR _0467_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[2\]
+ clknet_leaf_64_clk sg13g2_dfrbpq_2
X_5809_ VGND VPWR _2482_ _2486_ _0378_ _2487_ sg13g2_a21oi_1
XFILLER_11_926 VPWR VGND sg13g2_decap_8
XFILLER_10_436 VPWR VGND sg13g2_fill_1
X_6789_ net636 VGND VPWR _0398_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[6\]
+ clknet_leaf_58_clk sg13g2_dfrbpq_2
XFILLER_13_88 VPWR VGND sg13g2_fill_1
Xhold470 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[5\] VPWR
+ VGND net1227 sg13g2_dlygate4sd3_1
Xhold481 _1666_ VPWR VGND net1238 sg13g2_dlygate4sd3_1
Xhold492 _2580_ VPWR VGND net1249 sg13g2_dlygate4sd3_1
X_6658__64 VPWR VGND net64 sg13g2_tiehi
XFILLER_46_812 VPWR VGND sg13g2_fill_1
X_6399__380 VPWR VGND net564 sg13g2_tiehi
XFILLER_6_930 VPWR VGND sg13g2_decap_8
XFILLER_10_992 VPWR VGND sg13g2_decap_8
X_4140_ _1097_ VPWR _1105_ VGND net533 _0590_ sg13g2_o21ai_1
X_4071_ net445 _1055_ _0071_ VPWR VGND sg13g2_and2_1
XFILLER_49_672 VPWR VGND sg13g2_fill_2
XFILLER_48_182 VPWR VGND sg13g2_fill_2
XFILLER_37_856 VPWR VGND sg13g2_fill_2
X_4973_ _1798_ net1544 _1800_ VPWR VGND sg13g2_and2_1
X_3924_ net464 net825 _0054_ VPWR VGND sg13g2_and2_1
X_6712_ net713 VGND VPWR _0321_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[3\]
+ clknet_leaf_49_clk sg13g2_dfrbpq_1
X_6643_ net79 VGND VPWR _0252_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[4\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_1
X_3855_ _0885_ VPWR _0887_ VGND net1040 _0881_ sg13g2_o21ai_1
Xclkload9 clknet_4_12_0_clk clkload9/X VPWR VGND sg13g2_buf_8
X_6574_ net148 VGND VPWR net873 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[10\]
+ clknet_leaf_34_clk sg13g2_dfrbpq_2
X_3786_ _0833_ net929 net1056 VPWR VGND sg13g2_nand2b_1
X_5525_ _2245_ _2248_ _2249_ _2250_ VPWR VGND sg13g2_or3_1
X_5456_ VGND VPWR _2186_ _2190_ _2193_ _2189_ sg13g2_a21oi_1
X_4407_ _1321_ VPWR _1327_ VGND net542 _0603_ sg13g2_o21ai_1
X_5387_ net478 VPWR _2135_ VGND _2131_ _2134_ sg13g2_o21ai_1
X_4338_ _1266_ _1264_ _1269_ _1271_ VPWR VGND sg13g2_a21o_1
X_4269_ _1212_ _1213_ _1214_ VPWR VGND sg13g2_nor2b_1
X_6655__67 VPWR VGND net67 sg13g2_tiehi
X_6008_ _0413_ net460 _2650_ net1069 VPWR VGND sg13g2_and3_1
XFILLER_15_539 VPWR VGND sg13g2_fill_2
XFILLER_3_955 VPWR VGND sg13g2_decap_8
XFILLER_2_421 VPWR VGND sg13g2_fill_1
XFILLER_49_40 VPWR VGND sg13g2_decap_8
XFILLER_18_399 VPWR VGND sg13g2_fill_1
XFILLER_33_369 VPWR VGND sg13g2_fill_2
X_3640_ _0693_ _0683_ _0692_ VPWR VGND sg13g2_xnor2_1
X_3571_ hsync_sig _0626_ _0629_ VPWR VGND sg13g2_nand2_1
X_6473__249 VPWR VGND net249 sg13g2_tiehi
X_6290_ VGND VPWR net402 _2882_ _0466_ _2886_ sg13g2_a21oi_1
X_5310_ net837 net529 _2069_ VPWR VGND sg13g2_xor2_1
X_5241_ _2015_ _0565_ net379 VPWR VGND sg13g2_xnor2_1
X_5172_ _1947_ _1948_ _1955_ VPWR VGND sg13g2_nor2_1
X_4123_ net1222 net533 _1091_ VPWR VGND sg13g2_xor2_1
Xinput2 ui_in[0] net2 VPWR VGND sg13g2_buf_1
X_4054_ _1045_ _1038_ _1040_ VPWR VGND sg13g2_nand2_1
XFILLER_37_653 VPWR VGND sg13g2_fill_2
X_4956_ _1782_ _1785_ _1779_ _1786_ VPWR VGND sg13g2_nand3_1
X_4887_ VPWR _1728_ _1727_ VGND sg13g2_inv_1
X_3907_ _0921_ net1001 _0924_ VPWR VGND sg13g2_xor2_1
X_3838_ VGND VPWR net554 net857 _0020_ _0874_ sg13g2_a21oi_1
XFILLER_20_553 VPWR VGND sg13g2_fill_1
X_6626_ net96 VGND VPWR _0235_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[11\]
+ clknet_leaf_27_clk sg13g2_dfrbpq_1
X_6557_ net165 VGND VPWR net1136 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[7\]
+ clknet_leaf_40_clk sg13g2_dfrbpq_1
X_3769_ net419 net792 _0007_ VPWR VGND sg13g2_nor2_1
X_5508_ _2232_ _2230_ _2234_ _2236_ VPWR VGND sg13g2_a21o_1
X_6488_ net234 VGND VPWR net1357 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[2\]
+ clknet_leaf_50_clk sg13g2_dfrbpq_1
X_5439_ VGND VPWR _2171_ _2175_ _2178_ _2174_ sg13g2_a21oi_1
XFILLER_0_969 VPWR VGND sg13g2_decap_8
XFILLER_43_634 VPWR VGND sg13g2_fill_2
X_6797__444 VPWR VGND net628 sg13g2_tiehi
XFILLER_35_53 VPWR VGND sg13g2_fill_1
XFILLER_35_86 VPWR VGND sg13g2_fill_1
XFILLER_3_752 VPWR VGND sg13g2_decap_8
X_6880__325 VPWR VGND net325 sg13g2_tiehi
XFILLER_20_1024 VPWR VGND sg13g2_decap_4
XFILLER_33_111 VPWR VGND sg13g2_fill_1
X_4810_ _0202_ net471 _1663_ _1664_ VPWR VGND sg13g2_and3_1
X_5790_ VGND VPWR net1128 _2471_ _0374_ _2472_ sg13g2_a21oi_1
XFILLER_33_166 VPWR VGND sg13g2_fill_2
X_4741_ VGND VPWR _1602_ _1605_ _0191_ _1606_ sg13g2_a21oi_1
XFILLER_15_892 VPWR VGND sg13g2_decap_8
X_4672_ _1548_ _1543_ _1545_ VPWR VGND sg13g2_nand2b_1
X_6411_ net358 VGND VPWR net858 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[0\] clknet_leaf_65_clk
+ sg13g2_dfrbpq_1
X_3623_ _0676_ _0669_ _0675_ VPWR VGND sg13g2_xnor2_1
X_3554_ VPWR _0624_ net1130 VGND sg13g2_inv_1
X_6342_ net378 VPWR _2905_ VGND net844 _2903_ sg13g2_o21ai_1
X_6273_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[0\].y_shr\[0\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[0\].y_shr\[11\]
+ _2874_ VPWR VGND sg13g2_nor2_1
X_3485_ _0555_ net1566 VPWR VGND sg13g2_inv_2
X_5224_ _2000_ net1538 _1999_ VPWR VGND sg13g2_xnor2_1
X_5155_ _1942_ _1940_ _1941_ VPWR VGND sg13g2_nand2_1
X_5086_ net450 net14 _0260_ VPWR VGND sg13g2_and2_1
X_4106_ VGND VPWR net799 _1075_ _1077_ _1074_ sg13g2_a21oi_1
X_6449__295 VPWR VGND net295 sg13g2_tiehi
X_4037_ _1026_ VPWR _0063_ VGND net373 _1030_ sg13g2_o21ai_1
X_5988_ _2636_ net513 net1051 VPWR VGND sg13g2_xnor2_1
X_4939_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].z_sign u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[10\]
+ _1771_ VPWR VGND sg13g2_nor2b_1
X_6609_ net113 VGND VPWR net1252 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[7\]
+ clknet_leaf_25_clk sg13g2_dfrbpq_2
XFILLER_0_766 VPWR VGND sg13g2_decap_8
X_6428__324 VPWR VGND net324 sg13g2_tiehi
XFILLER_46_52 VPWR VGND sg13g2_fill_1
XFILLER_44_998 VPWR VGND sg13g2_fill_1
XFILLER_30_114 VPWR VGND sg13g2_fill_1
XFILLER_8_811 VPWR VGND sg13g2_decap_4
XFILLER_7_321 VPWR VGND sg13g2_fill_2
XFILLER_8_888 VPWR VGND sg13g2_decap_8
XFILLER_39_715 VPWR VGND sg13g2_fill_2
X_5911_ _2575_ _0576_ _0578_ _2562_ VPWR VGND sg13g2_and3_1
XFILLER_19_494 VPWR VGND sg13g2_fill_1
X_6891_ net726 VGND VPWR _0500_ u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[11\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
X_5842_ VPWR _2517_ _2516_ VGND sg13g2_inv_1
X_5773_ _2459_ net461 _2458_ VPWR VGND sg13g2_nand2_1
X_4724_ _1584_ net538 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[10\]
+ _1592_ VPWR VGND sg13g2_mux2_1
X_4655_ VGND VPWR _1530_ _1532_ _0177_ _1534_ sg13g2_a21oi_1
X_4586_ net437 _1475_ net1135 _0166_ VPWR VGND sg13g2_nor3_1
Xhold800 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[10\] VPWR VGND net1557
+ sg13g2_dlygate4sd3_1
Xhold811 _1240_ VPWR VGND net1568 sg13g2_dlygate4sd3_1
X_3606_ _0654_ _0658_ _0659_ VPWR VGND sg13g2_nor2_1
X_6787__454 VPWR VGND net638 sg13g2_tiehi
X_3537_ VPWR _0607_ net1110 VGND sg13g2_inv_1
X_6325_ net466 net796 _0496_ VPWR VGND sg13g2_and2_1
X_6256_ _2859_ net402 net555 _2860_ VPWR VGND sg13g2_a21o_2
X_3468_ VPWR _0538_ net983 VGND sg13g2_inv_1
X_5207_ _1985_ _0570_ _1984_ VPWR VGND sg13g2_xnor2_1
X_6187_ _2805_ _2806_ _0437_ VPWR VGND sg13g2_nor2b_1
X_5138_ VPWR VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[5\] _1911_
+ _1918_ _1906_ _1927_ _1913_ sg13g2_a221oi_1
X_5069_ _1879_ _1878_ _0246_ VPWR VGND sg13g2_nor2b_1
XFILLER_26_965 VPWR VGND sg13g2_decap_8
X_6794__447 VPWR VGND net631 sg13g2_tiehi
XFILLER_5_814 VPWR VGND sg13g2_decap_8
XFILLER_17_976 VPWR VGND sg13g2_decap_8
XFILLER_31_423 VPWR VGND sg13g2_fill_1
Xhold107 _0041_ VPWR VGND net864 sg13g2_dlygate4sd3_1
X_4440_ _1354_ _1355_ _1349_ _1356_ VPWR VGND sg13g2_nand3_1
Xhold118 _0875_ VPWR VGND net875 sg13g2_dlygate4sd3_1
Xhold129 _0063_ VPWR VGND net886 sg13g2_dlygate4sd3_1
X_6110_ _2739_ net1076 _2738_ VPWR VGND sg13g2_nand2_1
X_4371_ net503 VPWR _1298_ VGND _1296_ _1297_ sg13g2_o21ai_1
X_6041_ _2680_ net1295 _2678_ VPWR VGND sg13g2_xnor2_1
X_6874_ net337 VGND VPWR _0483_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[6\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_41_209 VPWR VGND sg13g2_fill_1
X_5825_ net457 VPWR _2502_ VGND _2495_ _2501_ sg13g2_o21ai_1
XFILLER_23_957 VPWR VGND sg13g2_decap_8
X_5756_ net472 VPWR _2445_ VGND _2443_ _2444_ sg13g2_o21ai_1
X_5687_ net516 _2386_ _2387_ VPWR VGND sg13g2_nor2_1
X_6492__230 VPWR VGND net230 sg13g2_tiehi
X_4707_ VGND VPWR _0609_ _1549_ _1577_ net537 sg13g2_a21oi_1
X_4638_ VGND VPWR _1520_ _1519_ _1513_ sg13g2_or2_1
Xhold630 _0311_ VPWR VGND net1387 sg13g2_dlygate4sd3_1
X_4569_ _1463_ net503 _1462_ VPWR VGND sg13g2_nand2_1
Xhold663 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[5\] VPWR
+ VGND net1420 sg13g2_dlygate4sd3_1
Xhold641 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[6\]\[5\] VPWR VGND net1398
+ sg13g2_dlygate4sd3_1
Xhold652 _0274_ VPWR VGND net1409 sg13g2_dlygate4sd3_1
Xhold674 _0243_ VPWR VGND net1431 sg13g2_dlygate4sd3_1
X_6308_ net446 net775 _0482_ VPWR VGND sg13g2_and2_1
Xhold685 _1406_ VPWR VGND net1442 sg13g2_dlygate4sd3_1
Xhold696 _0136_ VPWR VGND net1453 sg13g2_dlygate4sd3_1
X_6239_ _2846_ _2847_ _0448_ VPWR VGND sg13g2_nor2b_1
XFILLER_18_729 VPWR VGND sg13g2_fill_1
XFILLER_14_913 VPWR VGND sg13g2_decap_8
XFILLER_13_445 VPWR VGND sg13g2_fill_2
XFILLER_41_787 VPWR VGND sg13g2_fill_1
XFILLER_5_666 VPWR VGND sg13g2_fill_2
XFILLER_1_861 VPWR VGND sg13g2_decap_8
XFILLER_48_320 VPWR VGND sg13g2_fill_2
XFILLER_0_360 VPWR VGND sg13g2_fill_2
XFILLER_36_526 VPWR VGND sg13g2_fill_2
X_3940_ net450 VPWR _0055_ VGND _0932_ _0941_ sg13g2_o21ai_1
XFILLER_16_272 VPWR VGND sg13g2_fill_2
X_6777__464 VPWR VGND net648 sg13g2_tiehi
X_3871_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[6\] u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[5\]
+ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[0\] _0897_ VPWR VGND sg13g2_nor3_1
XFILLER_17_1018 VPWR VGND sg13g2_decap_8
X_6590_ net132 VGND VPWR net1366 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[1\]
+ clknet_leaf_25_clk sg13g2_dfrbpq_1
X_5610_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[7\] _2313_
+ _2321_ VPWR VGND sg13g2_nor2b_1
X_5541_ _2263_ net525 net1171 VPWR VGND sg13g2_xnor2_1
X_5472_ VPWR _2207_ _2206_ VGND sg13g2_inv_1
X_4423_ VGND VPWR _1334_ _1339_ _0138_ _1341_ sg13g2_a21oi_1
X_4354_ net1192 net541 _1284_ VPWR VGND sg13g2_xor2_1
X_6784__457 VPWR VGND net641 sg13g2_tiehi
Xfanout439 net440 net439 VPWR VGND sg13g2_buf_8
Xfanout417 _0562_ net417 VPWR VGND sg13g2_buf_2
Xfanout428 net440 net428 VPWR VGND sg13g2_buf_8
Xfanout406 _0644_ net406 VPWR VGND sg13g2_buf_8
X_6024_ _2659_ _2664_ _2665_ VPWR VGND sg13g2_nor2_1
X_4285_ _1226_ net1106 _1228_ VPWR VGND sg13g2_xor2_1
X_6857_ net371 VGND VPWR _0466_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[1\]
+ clknet_leaf_64_clk sg13g2_dfrbpq_2
XFILLER_11_905 VPWR VGND sg13g2_decap_8
X_5808_ net457 VPWR _2487_ VGND _2482_ _2486_ sg13g2_o21ai_1
X_6788_ net637 VGND VPWR net1437 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[5\]
+ clknet_leaf_58_clk sg13g2_dfrbpq_2
X_5739_ _2431_ net517 net877 VPWR VGND sg13g2_xnor2_1
Xhold460 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[12\] VPWR VGND net1217
+ sg13g2_dlygate4sd3_1
Xhold471 _2030_ VPWR VGND net1228 sg13g2_dlygate4sd3_1
Xhold493 _0393_ VPWR VGND net1250 sg13g2_dlygate4sd3_1
XFILLER_2_669 VPWR VGND sg13g2_decap_8
Xhold482 _0203_ VPWR VGND net1239 sg13g2_dlygate4sd3_1
XFILLER_38_20 VPWR VGND sg13g2_fill_1
XFILLER_38_97 VPWR VGND sg13g2_fill_2
XFILLER_18_537 VPWR VGND sg13g2_fill_1
XFILLER_13_297 VPWR VGND sg13g2_fill_2
XFILLER_10_971 VPWR VGND sg13g2_decap_8
XFILLER_6_986 VPWR VGND sg13g2_decap_8
X_4070_ _1053_ net840 _1055_ VPWR VGND sg13g2_xor2_1
XFILLER_37_813 VPWR VGND sg13g2_fill_2
X_6482__240 VPWR VGND net240 sg13g2_tiehi
X_4972_ net397 VPWR _1799_ VGND net1543 net1573 sg13g2_o21ai_1
X_6711_ net714 VGND VPWR net1389 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[2\]
+ clknet_leaf_56_clk sg13g2_dfrbpq_2
X_3923_ net463 net795 _0053_ VPWR VGND sg13g2_and2_1
X_3854_ net1040 _0881_ _0886_ VPWR VGND sg13g2_and2_1
X_6642_ net80 VGND VPWR _0251_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[3\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_1
X_6573_ net149 VGND VPWR net1178 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[2\]
+ clknet_leaf_33_clk sg13g2_dfrbpq_2
X_3785_ _0832_ _0549_ net978 _0548_ net920 VPWR VGND sg13g2_a22oi_1
X_5524_ _2243_ _2244_ _2249_ VPWR VGND sg13g2_nor2_1
X_5455_ _2191_ _2192_ _0319_ VPWR VGND sg13g2_and2_1
X_4406_ _1324_ _1320_ _1323_ _1326_ VPWR VGND sg13g2_a21o_1
X_5386_ _2132_ net1390 _2134_ VPWR VGND sg13g2_xor2_1
X_4337_ _1266_ _1269_ _1264_ _1270_ VPWR VGND sg13g2_nand3_1
X_4268_ VGND VPWR _1213_ _1211_ net1501 sg13g2_or2_1
X_6007_ net414 VPWR _2651_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[9\]
+ net1068 sg13g2_o21ai_1
X_4199_ _1155_ net991 _1154_ VPWR VGND sg13g2_nand2_1
XFILLER_28_846 VPWR VGND sg13g2_fill_2
XFILLER_39_194 VPWR VGND sg13g2_fill_1
XFILLER_43_816 VPWR VGND sg13g2_fill_1
X_6598__124 VPWR VGND net124 sg13g2_tiehi
XFILLER_42_348 VPWR VGND sg13g2_fill_1
X_6909_ net282 VGND VPWR _0504_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[3\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_23_562 VPWR VGND sg13g2_fill_1
XFILLER_7_706 VPWR VGND sg13g2_fill_2
X_6459__275 VPWR VGND net275 sg13g2_tiehi
XFILLER_3_934 VPWR VGND sg13g2_decap_8
XFILLER_2_466 VPWR VGND sg13g2_fill_1
X_6767__474 VPWR VGND net658 sg13g2_tiehi
Xhold290 _2653_ VPWR VGND net1047 sg13g2_dlygate4sd3_1
XFILLER_49_96 VPWR VGND sg13g2_fill_2
XFILLER_34_827 VPWR VGND sg13g2_fill_2
X_6698__557 VPWR VGND net741 sg13g2_tiehi
X_6774__467 VPWR VGND net651 sg13g2_tiehi
XFILLER_41_381 VPWR VGND sg13g2_fill_2
X_3570_ u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[8\] _0541_ _0627_ _0628_ _0629_ VPWR
+ VGND sg13g2_nor4_1
XFILLER_6_783 VPWR VGND sg13g2_decap_8
XFILLER_5_271 VPWR VGND sg13g2_fill_1
X_5240_ _2014_ net1181 net379 VPWR VGND sg13g2_nand2_1
X_5171_ VGND VPWR _1952_ _1953_ _0273_ _1954_ sg13g2_a21oi_1
X_4122_ VGND VPWR _1086_ _1088_ _0088_ _1090_ sg13g2_a21oi_1
X_4053_ _1044_ net982 net376 VPWR VGND sg13g2_nand2_1
Xinput3 ui_in[1] net3 VPWR VGND sg13g2_buf_1
XFILLER_37_621 VPWR VGND sg13g2_fill_1
X_6896__547 VPWR VGND net731 sg13g2_tiehi
X_4955_ _1785_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[3\] net399
+ VPWR VGND sg13g2_xnor2_1
X_3906_ _0923_ net1001 _0885_ VPWR VGND sg13g2_nand2_1
X_4886_ net389 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[5\] _1727_
+ VPWR VGND sg13g2_xor2_1
X_3837_ net441 VPWR _0874_ VGND net554 net857 sg13g2_o21ai_1
X_6625_ net97 VGND VPWR _0234_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[10\]
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
X_6556_ net166 VGND VPWR _0165_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[6\]
+ clknet_leaf_39_clk sg13g2_dfrbpq_1
X_3768_ net553 net813 _0006_ VPWR VGND sg13g2_nor2b_1
X_5507_ _2232_ _2234_ _2230_ _2235_ VPWR VGND sg13g2_nand3_1
X_6487_ net235 VGND VPWR net1105 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[1\]
+ clknet_leaf_51_clk sg13g2_dfrbpq_2
X_3699_ VPWR _0752_ _0751_ VGND sg13g2_inv_1
X_5438_ _2176_ _2177_ _0317_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_948 VPWR VGND sg13g2_decap_8
X_5369_ net522 _2118_ _2119_ VPWR VGND sg13g2_nor2_1
XFILLER_19_77 VPWR VGND sg13g2_fill_1
X_6651__71 VPWR VGND net71 sg13g2_tiehi
XFILLER_23_381 VPWR VGND sg13g2_fill_1
XFILLER_13_1021 VPWR VGND sg13g2_decap_8
XFILLER_3_731 VPWR VGND sg13g2_decap_8
XFILLER_39_919 VPWR VGND sg13g2_fill_1
XFILLER_20_1003 VPWR VGND sg13g2_decap_8
XFILLER_18_186 VPWR VGND sg13g2_fill_2
X_4740_ net488 VPWR _1606_ VGND _1602_ _1605_ sg13g2_o21ai_1
X_4671_ _1547_ net1534 net393 VPWR VGND sg13g2_xnor2_1
X_6410_ net360 VGND VPWR net891 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[8\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
X_3622_ _0673_ _0657_ _0675_ VPWR VGND sg13g2_xor2_1
X_6341_ net374 _2903_ net927 _0505_ VPWR VGND sg13g2_nor3_1
X_3553_ VPWR _0623_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[9\] VGND
+ sg13g2_inv_1
XFILLER_44_0 VPWR VGND sg13g2_fill_1
X_6272_ _2867_ _2872_ _2873_ VPWR VGND sg13g2_nor2_2
X_3484_ VPWR _0554_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[1\] VGND
+ sg13g2_inv_1
X_5223_ _1999_ _1998_ _1997_ VPWR VGND sg13g2_nand2b_1
X_6588__134 VPWR VGND net134 sg13g2_tiehi
X_5154_ _1941_ net1558 net380 VPWR VGND sg13g2_xnor2_1
X_4105_ VGND VPWR net799 _1075_ _0085_ _1076_ sg13g2_a21oi_1
X_5085_ net450 net13 _0259_ VPWR VGND sg13g2_and2_1
X_4036_ _1030_ _1027_ _1029_ VPWR VGND sg13g2_xnor2_1
XFILLER_13_808 VPWR VGND sg13g2_fill_1
X_5987_ _2635_ net513 net1051 VPWR VGND sg13g2_nand2_1
X_4938_ net426 net947 _0224_ VPWR VGND sg13g2_nor2_1
X_6595__127 VPWR VGND net127 sg13g2_tiehi
X_4869_ _1713_ _1712_ _1709_ VPWR VGND sg13g2_nand2b_1
X_6757__484 VPWR VGND net668 sg13g2_tiehi
X_6608_ net114 VGND VPWR _0217_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[6\]
+ clknet_leaf_24_clk sg13g2_dfrbpq_1
XFILLER_4_528 VPWR VGND sg13g2_fill_2
X_6539_ net183 VGND VPWR net1226 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[2\]
+ clknet_leaf_33_clk sg13g2_dfrbpq_1
X_6688__567 VPWR VGND net751 sg13g2_tiehi
XFILLER_0_745 VPWR VGND sg13g2_decap_8
X_6764__477 VPWR VGND net661 sg13g2_tiehi
XFILLER_48_738 VPWR VGND sg13g2_fill_2
XFILLER_8_867 VPWR VGND sg13g2_decap_8
XFILLER_39_705 VPWR VGND sg13g2_fill_1
XFILLER_38_215 VPWR VGND sg13g2_fill_1
XFILLER_38_226 VPWR VGND sg13g2_fill_1
XFILLER_47_760 VPWR VGND sg13g2_fill_1
X_5910_ VGND VPWR _2568_ _2572_ _2574_ _2571_ sg13g2_a21oi_1
X_6890_ net292 VGND VPWR _0499_ u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[10\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
X_5841_ _2516_ net1306 _2514_ VPWR VGND sg13g2_xnor2_1
XFILLER_22_627 VPWR VGND sg13g2_fill_2
X_5772_ VGND VPWR _2458_ _2457_ _2455_ sg13g2_or2_1
XFILLER_34_498 VPWR VGND sg13g2_fill_2
X_4723_ _1591_ _1586_ _1590_ VPWR VGND sg13g2_nand2_1
X_4654_ _1534_ net481 _1533_ VPWR VGND sg13g2_nand2_1
Xhold812 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[12\] VPWR VGND net1569
+ sg13g2_dlygate4sd3_1
X_4585_ VGND VPWR _1470_ _1472_ _1476_ net1134 sg13g2_a21oi_1
Xhold801 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[8\] VPWR VGND net1558
+ sg13g2_dlygate4sd3_1
X_3605_ _0658_ _0638_ _0656_ VPWR VGND sg13g2_xnor2_1
X_6324_ net462 net771 _0495_ VPWR VGND sg13g2_and2_1
X_3536_ VPWR _0606_ net1120 VGND sg13g2_inv_1
X_6255_ _2859_ net967 _0605_ VPWR VGND sg13g2_nand2_1
XFILLER_27_1009 VPWR VGND sg13g2_decap_8
X_3467_ VPWR _0537_ net1024 VGND sg13g2_inv_1
X_5206_ VGND VPWR net415 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[8\]
+ _1984_ _1977_ sg13g2_a21oi_1
X_6186_ VGND VPWR _2800_ _2804_ _2806_ net424 sg13g2_a21oi_1
X_5137_ _1926_ net1162 _1925_ VPWR VGND sg13g2_xnor2_1
X_5068_ net464 VPWR _1879_ VGND _1876_ _1877_ sg13g2_o21ai_1
X_4019_ _1015_ net961 net377 VPWR VGND sg13g2_nand2_1
XFILLER_13_616 VPWR VGND sg13g2_fill_2
X_6462__271 VPWR VGND net271 sg13g2_tiehi
XFILLER_32_66 VPWR VGND sg13g2_fill_2
XFILLER_10_1013 VPWR VGND sg13g2_decap_8
XFILLER_0_520 VPWR VGND sg13g2_fill_2
XFILLER_17_955 VPWR VGND sg13g2_decap_8
X_6578__144 VPWR VGND net144 sg13g2_tiehi
X_6916__266 VPWR VGND net266 sg13g2_tiehi
XFILLER_8_697 VPWR VGND sg13g2_fill_2
Xhold108 u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[9\] VPWR VGND net865 sg13g2_dlygate4sd3_1
Xhold119 _0021_ VPWR VGND net876 sg13g2_dlygate4sd3_1
X_4370_ _1297_ net541 net1121 VPWR VGND sg13g2_xnor2_1
XFILLER_4_881 VPWR VGND sg13g2_decap_8
X_6585__137 VPWR VGND net137 sg13g2_tiehi
X_6040_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[4\] _2678_ _2679_
+ VPWR VGND sg13g2_and2_1
XFILLER_3_391 VPWR VGND sg13g2_fill_1
X_6747__494 VPWR VGND net678 sg13g2_tiehi
XFILLER_39_513 VPWR VGND sg13g2_fill_2
XFILLER_35_730 VPWR VGND sg13g2_fill_1
X_6873_ net339 VGND VPWR _0482_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[5\]
+ clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5824_ _2501_ net1348 _2499_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_936 VPWR VGND sg13g2_decap_8
XFILLER_35_796 VPWR VGND sg13g2_fill_1
XFILLER_31_991 VPWR VGND sg13g2_fill_1
X_5755_ _2439_ VPWR _2444_ VGND _2437_ _2438_ sg13g2_o21ai_1
X_4706_ VGND VPWR _1569_ _1573_ _1576_ _1572_ sg13g2_a21oi_1
X_5686_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[8\] _2373_ _2386_
+ VPWR VGND sg13g2_nor2_1
X_6754__487 VPWR VGND net671 sg13g2_tiehi
XFILLER_30_490 VPWR VGND sg13g2_fill_2
X_4637_ _1519_ net1212 _1517_ VPWR VGND sg13g2_xnor2_1
Xhold620 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[2\] VPWR
+ VGND net1377 sg13g2_dlygate4sd3_1
Xhold642 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[12\] VPWR VGND net1399
+ sg13g2_dlygate4sd3_1
Xhold653 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[7\] VPWR VGND net1410
+ sg13g2_dlygate4sd3_1
Xhold631 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[3\] VPWR
+ VGND net1388 sg13g2_dlygate4sd3_1
X_4568_ VGND VPWR _1462_ _1461_ _1460_ sg13g2_or2_1
Xhold675 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[6\] VPWR VGND net1432
+ sg13g2_dlygate4sd3_1
Xhold697 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[4\] VPWR
+ VGND net1454 sg13g2_dlygate4sd3_1
Xhold686 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[1\] VPWR
+ VGND net1443 sg13g2_dlygate4sd3_1
X_4499_ _1406_ _0602_ _1404_ VPWR VGND sg13g2_nand2_1
X_6307_ net454 net786 _0481_ VPWR VGND sg13g2_and2_1
X_3519_ VPWR _0589_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[6\] VGND
+ sg13g2_inv_1
Xhold664 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[8\] VPWR VGND net1421
+ sg13g2_dlygate4sd3_1
X_6238_ VGND VPWR _2844_ _2845_ _2847_ net424 sg13g2_a21oi_1
X_6169_ _2786_ _2790_ _2791_ VPWR VGND sg13g2_nor2_1
XFILLER_14_969 VPWR VGND sg13g2_decap_8
XFILLER_40_265 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_20_clk clknet_4_5_0_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
XFILLER_5_623 VPWR VGND sg13g2_fill_1
XFILLER_4_155 VPWR VGND sg13g2_fill_1
XFILLER_1_840 VPWR VGND sg13g2_decap_8
XFILLER_1_1022 VPWR VGND sg13g2_decap_8
X_3870_ VGND VPWR _0538_ _0894_ _0030_ _0896_ sg13g2_a21oi_1
X_5540_ net525 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[9\] _2262_
+ VPWR VGND sg13g2_nor2b_1
Xclkbuf_leaf_11_clk clknet_4_6_0_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
XFILLER_9_995 VPWR VGND sg13g2_decap_8
X_5471_ _2200_ net522 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[12\]
+ _2206_ VPWR VGND sg13g2_mux2_1
X_4422_ _1341_ net496 _1340_ VPWR VGND sg13g2_nand2_1
X_4353_ _1283_ net410 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[6\]
+ VPWR VGND sg13g2_nand2_1
X_6667__55 VPWR VGND net55 sg13g2_tiehi
X_4284_ _1226_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[6\] _1227_
+ VPWR VGND sg13g2_nor2b_1
Xfanout418 _0553_ net418 VPWR VGND sg13g2_buf_8
Xfanout429 net434 net429 VPWR VGND sg13g2_buf_8
Xfanout407 _0643_ net407 VPWR VGND sg13g2_buf_8
X_6023_ _2662_ _2663_ _2664_ VPWR VGND sg13g2_nor2b_1
X_6856_ net557 VGND VPWR _0465_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[0\]
+ clknet_leaf_64_clk sg13g2_dfrbpq_2
X_3999_ _0993_ VPWR _0057_ VGND _0996_ _0998_ sg13g2_o21ai_1
X_5807_ _2486_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[2\] _2484_
+ VPWR VGND sg13g2_xnor2_1
X_6787_ net638 VGND VPWR net1555 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[4\]
+ clknet_leaf_58_clk sg13g2_dfrbpq_1
XFILLER_13_57 VPWR VGND sg13g2_fill_1
X_5738_ net517 net877 _2430_ VPWR VGND sg13g2_nor2b_1
X_5669_ _2367_ VPWR _2371_ VGND _2364_ _2369_ sg13g2_o21ai_1
Xhold450 _0149_ VPWR VGND net1207 sg13g2_dlygate4sd3_1
Xhold461 _0388_ VPWR VGND net1218 sg13g2_dlygate4sd3_1
Xhold472 _0286_ VPWR VGND net1229 sg13g2_dlygate4sd3_1
Xhold494 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[6\] VPWR VGND net1251
+ sg13g2_dlygate4sd3_1
Xhold483 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[3\]\[1\] VPWR VGND net1240
+ sg13g2_dlygate4sd3_1
X_6568__154 VPWR VGND net154 sg13g2_tiehi
X_6575__147 VPWR VGND net147 sg13g2_tiehi
XFILLER_10_950 VPWR VGND sg13g2_decap_8
XFILLER_6_965 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
X_6664__58 VPWR VGND net58 sg13g2_tiehi
XFILLER_49_674 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_0_clk clknet_4_0_0_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
X_6744__497 VPWR VGND net681 sg13g2_tiehi
X_4971_ _1798_ _1792_ _1796_ VPWR VGND sg13g2_nand2_1
X_3922_ net463 net788 _0052_ VPWR VGND sg13g2_and2_1
X_6710_ net715 VGND VPWR _0319_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[1\]
+ clknet_leaf_55_clk sg13g2_dfrbpq_2
X_3853_ net419 _0884_ _0885_ VPWR VGND sg13g2_nor2_2
X_6641_ net81 VGND VPWR _0250_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[2\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_1
X_6790__451 VPWR VGND net635 sg13g2_tiehi
X_3784_ _0831_ net944 net1003 VPWR VGND sg13g2_nand2b_1
X_6572_ net150 VGND VPWR _0181_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[1\]
+ clknet_leaf_33_clk sg13g2_dfrbpq_2
X_5523_ _2248_ net523 net1506 VPWR VGND sg13g2_xnor2_1
XFILLER_30_1027 VPWR VGND sg13g2_fill_2
X_5454_ VGND VPWR _2186_ _2190_ _2192_ net429 sg13g2_a21oi_1
X_5385_ net1390 _2132_ _2133_ VPWR VGND sg13g2_nor2_1
X_4405_ VGND VPWR _1320_ _1324_ _0136_ _1325_ sg13g2_a21oi_1
X_4336_ net1284 net542 _1269_ VPWR VGND sg13g2_xor2_1
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
X_4267_ net1501 _1211_ _1212_ VPWR VGND sg13g2_and2_1
X_6006_ _2650_ _2648_ _2645_ VPWR VGND sg13g2_nand2b_1
X_4198_ _1154_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[12\] _1152_
+ VPWR VGND sg13g2_xnor2_1
X_6908_ net284 VGND VPWR net900 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[2\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_1
X_6839_ net586 VGND VPWR _0448_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[8\]
+ clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_10_202 VPWR VGND sg13g2_fill_2
XFILLER_11_747 VPWR VGND sg13g2_fill_1
XFILLER_3_913 VPWR VGND sg13g2_decap_8
Xhold280 _1114_ VPWR VGND net1037 sg13g2_dlygate4sd3_1
Xhold291 _0414_ VPWR VGND net1048 sg13g2_dlygate4sd3_1
XFILLER_49_75 VPWR VGND sg13g2_decap_8
XFILLER_6_762 VPWR VGND sg13g2_decap_8
XFILLER_5_250 VPWR VGND sg13g2_fill_1
X_5170_ net493 VPWR _1954_ VGND _1952_ _1953_ sg13g2_o21ai_1
X_4121_ _1090_ net501 _1089_ VPWR VGND sg13g2_nand2_1
X_4052_ net376 net1012 _1043_ _0065_ VPWR VGND sg13g2_a21o_1
Xinput4 ui_in[2] net4 VPWR VGND sg13g2_buf_1
X_4954_ VGND VPWR _1784_ net399 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[3\]
+ sg13g2_or2_1
X_3905_ net420 net915 _0922_ _0039_ VPWR VGND sg13g2_nor3_1
X_4885_ VGND VPWR net1167 net389 _1726_ _1724_ sg13g2_a21oi_1
X_6558__164 VPWR VGND net164 sg13g2_tiehi
X_3836_ net890 VPWR _0019_ VGND _0870_ _0873_ sg13g2_o21ai_1
X_6624_ net98 VGND VPWR net1187 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[9\]
+ clknet_leaf_27_clk sg13g2_dfrbpq_1
X_6555_ net167 VGND VPWR _0164_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[5\]
+ clknet_leaf_40_clk sg13g2_dfrbpq_1
X_3767_ net553 net835 _0005_ VPWR VGND sg13g2_nor2b_1
X_5506_ _2234_ net524 net1089 VPWR VGND sg13g2_xnor2_1
X_6486_ net236 VGND VPWR _0095_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[0\]
+ clknet_leaf_36_clk sg13g2_dfrbpq_1
XFILLER_10_36 VPWR VGND sg13g2_fill_2
X_3698_ _0686_ net403 _0751_ VPWR VGND sg13g2_xor2_1
X_5437_ VGND VPWR _2171_ _2175_ _2177_ net429 sg13g2_a21oi_1
XFILLER_0_927 VPWR VGND sg13g2_decap_8
X_5368_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[5\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[6\]
+ _2095_ _2118_ VPWR VGND sg13g2_nor3_1
X_4319_ _1234_ VPWR _1256_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[10\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[11\] sg13g2_o21ai_1
X_5299_ net1313 net529 _2060_ VPWR VGND sg13g2_xor2_1
X_6565__157 VPWR VGND net157 sg13g2_tiehi
XFILLER_13_1000 VPWR VGND sg13g2_decap_8
X_6396__385 VPWR VGND net569 sg13g2_tiehi
XFILLER_3_710 VPWR VGND sg13g2_decap_8
X_6472__251 VPWR VGND net251 sg13g2_tiehi
XFILLER_3_787 VPWR VGND sg13g2_decap_8
X_6780__461 VPWR VGND net645 sg13g2_tiehi
XFILLER_46_496 VPWR VGND sg13g2_fill_1
XFILLER_33_168 VPWR VGND sg13g2_fill_1
XFILLER_30_864 VPWR VGND sg13g2_fill_1
X_4670_ VGND VPWR _1544_ _1545_ _0180_ _1546_ sg13g2_a21oi_1
X_3621_ _0657_ _0673_ _0674_ VPWR VGND sg13g2_nor2_1
X_3552_ VPWR _0622_ net1536 VGND sg13g2_inv_1
X_6340_ net926 _2901_ _2904_ VPWR VGND sg13g2_nor2_1
X_6271_ _2870_ _2871_ _2872_ VPWR VGND sg13g2_and2_1
X_3483_ _0553_ net523 VPWR VGND sg13g2_inv_2
X_5222_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[11\] VPWR _1998_ VGND
+ _1991_ _1996_ sg13g2_o21ai_1
X_5153_ _1938_ _1931_ _1937_ _1940_ VPWR VGND sg13g2_a21o_1
XFILLER_37_0 VPWR VGND sg13g2_fill_2
X_4104_ net499 VPWR _1076_ VGND net799 _1075_ sg13g2_o21ai_1
X_5084_ net449 net12 _0258_ VPWR VGND sg13g2_and2_1
XFILLER_37_452 VPWR VGND sg13g2_fill_2
X_4035_ _1029_ _0937_ _1028_ VPWR VGND sg13g2_nand2_1
X_5986_ VGND VPWR net810 _2632_ _2634_ _2631_ sg13g2_a21oi_1
X_4937_ _1770_ net946 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[10\]
+ VPWR VGND sg13g2_xnor2_1
X_4868_ _1712_ _0616_ _1711_ VPWR VGND sg13g2_xnor2_1
X_6607_ net115 VGND VPWR net1168 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[5\]
+ clknet_leaf_24_clk sg13g2_dfrbpq_1
XFILLER_20_374 VPWR VGND sg13g2_fill_2
X_3819_ _0859_ _0807_ _0814_ VPWR VGND sg13g2_nand2_1
X_4799_ _1653_ _1654_ _1655_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_396 VPWR VGND sg13g2_fill_2
X_6538_ net184 VGND VPWR net997 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[1\]
+ clknet_leaf_32_clk sg13g2_dfrbpq_1
X_6469_ net257 VGND VPWR _0078_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[8\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_0_724 VPWR VGND sg13g2_decap_8
XFILLER_48_728 VPWR VGND sg13g2_fill_1
XFILLER_46_10 VPWR VGND sg13g2_fill_1
XFILLER_29_997 VPWR VGND sg13g2_decap_8
XFILLER_31_628 VPWR VGND sg13g2_fill_2
XFILLER_8_846 VPWR VGND sg13g2_decap_8
XFILLER_7_323 VPWR VGND sg13g2_fill_1
XFILLER_12_886 VPWR VGND sg13g2_decap_8
XFILLER_39_717 VPWR VGND sg13g2_fill_1
X_6548__174 VPWR VGND net174 sg13g2_tiehi
XFILLER_35_956 VPWR VGND sg13g2_fill_2
XFILLER_35_967 VPWR VGND sg13g2_fill_2
X_5840_ net1306 _2514_ _2515_ VPWR VGND sg13g2_and2_1
X_5771_ net1078 net518 _2457_ VPWR VGND sg13g2_xor2_1
X_4722_ _0188_ net488 _1589_ _1590_ VPWR VGND sg13g2_and3_1
X_6856__373 VPWR VGND net557 sg13g2_tiehi
X_6555__167 VPWR VGND net167 sg13g2_tiehi
X_4653_ VGND VPWR _1533_ _1532_ _1530_ sg13g2_or2_1
Xhold802 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[3\] VPWR
+ VGND net1559 sg13g2_dlygate4sd3_1
X_3604_ _0657_ _0638_ _0656_ VPWR VGND sg13g2_nand2_1
X_4584_ _1475_ _1470_ _1472_ _1474_ VPWR VGND sg13g2_and3_1
X_6323_ net468 net801 _0494_ VPWR VGND sg13g2_and2_1
X_3535_ VPWR _0605_ net506 VGND sg13g2_inv_1
XFILLER_7_890 VPWR VGND sg13g2_decap_8
Xhold813 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[9\] VPWR VGND net1570
+ sg13g2_dlygate4sd3_1
X_6254_ VGND VPWR net402 net968 _0452_ net421 sg13g2_a21oi_1
X_3466_ VPWR _0536_ net920 VGND sg13g2_inv_1
X_5205_ _1979_ VPWR _1983_ VGND _1976_ _1981_ sg13g2_o21ai_1
X_6185_ _2800_ _2804_ _2805_ VPWR VGND sg13g2_nor2_1
X_5136_ _1923_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[6\]
+ _1925_ VPWR VGND sg13g2_xor2_1
X_5067_ _1878_ _1876_ _1877_ VPWR VGND sg13g2_nand2_1
X_4018_ _1010_ VPWR _0060_ VGND net372 _1014_ sg13g2_o21ai_1
XFILLER_26_956 VPWR VGND sg13g2_fill_1
X_5969_ VGND VPWR _2617_ _2621_ _2626_ _2624_ sg13g2_a21oi_1
X_6694__561 VPWR VGND net745 sg13g2_tiehi
XFILLER_32_34 VPWR VGND sg13g2_fill_2
X_6770__471 VPWR VGND net655 sg13g2_tiehi
XFILLER_5_849 VPWR VGND sg13g2_decap_8
XFILLER_17_934 VPWR VGND sg13g2_decap_8
X_6886__300 VPWR VGND net300 sg13g2_tiehi
Xhold109 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[6\] VPWR VGND net866 sg13g2_dlygate4sd3_1
XFILLER_4_860 VPWR VGND sg13g2_decap_8
XFILLER_26_1021 VPWR VGND sg13g2_decap_8
XFILLER_39_569 VPWR VGND sg13g2_fill_1
XFILLER_35_720 VPWR VGND sg13g2_fill_1
X_6872_ net341 VGND VPWR _0481_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[4\]
+ clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5823_ _2500_ net1348 _2499_ VPWR VGND sg13g2_nand2_1
XFILLER_22_403 VPWR VGND sg13g2_fill_2
X_5754_ _2443_ net517 net1204 VPWR VGND sg13g2_xnor2_1
X_4705_ net1439 _1575_ _0186_ VPWR VGND sg13g2_nor2b_1
X_5685_ _2382_ VPWR _2385_ VGND _2379_ _2383_ sg13g2_o21ai_1
X_4636_ _1518_ net1212 _1517_ VPWR VGND sg13g2_nand2_2
Xhold621 _0356_ VPWR VGND net1378 sg13g2_dlygate4sd3_1
Xhold610 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[4\]\[3\] VPWR VGND net1367
+ sg13g2_dlygate4sd3_1
Xhold643 _0196_ VPWR VGND net1400 sg13g2_dlygate4sd3_1
X_4567_ _1456_ VPWR _1461_ VGND _1454_ _1455_ sg13g2_o21ai_1
Xhold632 _0320_ VPWR VGND net1389 sg13g2_dlygate4sd3_1
X_6306_ net462 net769 _0480_ VPWR VGND sg13g2_and2_1
Xhold654 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[5\] VPWR VGND net1411
+ sg13g2_dlygate4sd3_1
Xhold687 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[7\] VPWR VGND net1444
+ sg13g2_dlygate4sd3_1
XFILLER_1_318 VPWR VGND sg13g2_fill_2
XFILLER_1_329 VPWR VGND sg13g2_fill_1
Xhold665 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[10\] VPWR VGND net1422
+ sg13g2_dlygate4sd3_1
X_3518_ VPWR _0588_ net1154 VGND sg13g2_inv_1
Xhold676 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[7\] VPWR VGND net1433
+ sg13g2_dlygate4sd3_1
X_4498_ _0602_ _1404_ _1405_ VPWR VGND sg13g2_nor2_1
Xhold698 _2593_ VPWR VGND net1455 sg13g2_dlygate4sd3_1
X_6237_ _2844_ _2845_ _2846_ VPWR VGND sg13g2_nor2_1
X_6168_ _2790_ _0622_ _2788_ VPWR VGND sg13g2_xnor2_1
X_5119_ _1910_ net1275 _1909_ VPWR VGND sg13g2_nand2_1
X_6099_ _2728_ _2730_ _0425_ VPWR VGND sg13g2_nor2_1
XFILLER_14_948 VPWR VGND sg13g2_decap_8
XFILLER_43_99 VPWR VGND sg13g2_fill_2
XFILLER_43_66 VPWR VGND sg13g2_fill_2
X_6538__184 VPWR VGND net184 sg13g2_tiehi
XFILLER_49_1021 VPWR VGND sg13g2_decap_8
XFILLER_5_668 VPWR VGND sg13g2_fill_1
XFILLER_1_896 VPWR VGND sg13g2_decap_8
X_6545__177 VPWR VGND net177 sg13g2_tiehi
XFILLER_1_1001 VPWR VGND sg13g2_decap_8
X_6591__131 VPWR VGND net131 sg13g2_tiehi
XFILLER_9_974 VPWR VGND sg13g2_decap_8
X_5470_ _0321_ net479 _2204_ _2205_ VPWR VGND sg13g2_and3_1
X_4421_ VGND VPWR _1340_ _1339_ _1334_ sg13g2_or2_1
X_4352_ _1280_ _1281_ _1282_ VPWR VGND sg13g2_nor2_1
Xfanout419 net423 net419 VPWR VGND sg13g2_buf_8
X_4283_ _1226_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[10\]
+ _1224_ VPWR VGND sg13g2_xnor2_1
Xfanout408 _0642_ net408 VPWR VGND sg13g2_buf_8
X_6022_ VGND VPWR _2663_ _2661_ net1264 sg13g2_or2_1
X_6684__571 VPWR VGND net755 sg13g2_tiehi
X_6760__481 VPWR VGND net665 sg13g2_tiehi
X_6855_ net560 VGND VPWR _0464_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[12\]
+ clknet_leaf_7_clk sg13g2_dfrbpq_2
X_3998_ _0992_ VPWR _0998_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[0\]
+ _0995_ sg13g2_o21ai_1
X_5806_ _2485_ net1474 _2484_ VPWR VGND sg13g2_nand2_1
X_6786_ net639 VGND VPWR _0395_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[3\]
+ clknet_leaf_60_clk sg13g2_dfrbpq_2
X_5737_ net809 net427 _0364_ VPWR VGND sg13g2_nor2_1
X_6691__564 VPWR VGND net748 sg13g2_tiehi
X_5668_ VGND VPWR _2364_ _2369_ _0354_ _2370_ sg13g2_a21oi_1
X_4619_ _1501_ net1382 _1503_ VPWR VGND sg13g2_xor2_1
X_5599_ VGND VPWR _2306_ net1413 _0344_ _2311_ sg13g2_a21oi_1
Xhold462 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[8\] VPWR VGND net1219
+ sg13g2_dlygate4sd3_1
Xhold440 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[11\] VPWR VGND net1197
+ sg13g2_dlygate4sd3_1
Xhold451 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[1\] VPWR
+ VGND net1208 sg13g2_dlygate4sd3_1
Xhold495 _0218_ VPWR VGND net1252 sg13g2_dlygate4sd3_1
Xhold473 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[0\] VPWR
+ VGND net1230 sg13g2_dlygate4sd3_1
Xhold484 _0352_ VPWR VGND net1241 sg13g2_dlygate4sd3_1
X_6906__288 VPWR VGND net288 sg13g2_tiehi
XFILLER_14_734 VPWR VGND sg13g2_fill_1
XFILLER_6_944 VPWR VGND sg13g2_decap_8
XFILLER_49_620 VPWR VGND sg13g2_fill_2
XFILLER_1_693 VPWR VGND sg13g2_decap_8
XFILLER_23_1013 VPWR VGND sg13g2_decap_8
XFILLER_36_358 VPWR VGND sg13g2_fill_1
X_4970_ VGND VPWR _1794_ _1795_ _0229_ _1797_ sg13g2_a21oi_1
X_3921_ net465 net807 _0051_ VPWR VGND sg13g2_and2_1
X_3852_ _0884_ _0827_ _0881_ _0883_ VPWR VGND sg13g2_and3_2
X_6640_ net82 VGND VPWR _0249_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[1\]
+ clknet_leaf_14_clk sg13g2_dfrbpq_2
X_6571_ net151 VGND VPWR _0180_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[0\]
+ clknet_leaf_33_clk sg13g2_dfrbpq_2
X_3783_ net554 net1065 _0830_ VPWR VGND sg13g2_nor2b_1
XFILLER_30_1006 VPWR VGND sg13g2_decap_8
X_5522_ VGND VPWR _2243_ _2246_ _0331_ _2247_ sg13g2_a21oi_1
X_5453_ VGND VPWR _2191_ _2190_ _2186_ sg13g2_or2_1
X_5384_ _2125_ net522 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[10\]
+ _2132_ VPWR VGND sg13g2_mux2_1
X_4404_ net497 VPWR _1325_ VGND _1320_ _1324_ sg13g2_o21ai_1
X_4335_ _1268_ net410 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[3\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_8_1007 VPWR VGND sg13g2_decap_8
X_4266_ _1211_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[4\]
+ _1209_ VPWR VGND sg13g2_xnor2_1
X_6005_ VGND VPWR _2647_ _2648_ _0412_ _2649_ sg13g2_a21oi_1
X_4197_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[12\] _1152_ _1153_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_28_848 VPWR VGND sg13g2_fill_1
X_6528__194 VPWR VGND net194 sg13g2_tiehi
X_6907_ net286 VGND VPWR _0502_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[1\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_1
XFILLER_36_892 VPWR VGND sg13g2_fill_2
X_6838_ net587 VGND VPWR _0447_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[7\]
+ clknet_leaf_11_clk sg13g2_dfrbpq_1
X_6769_ net656 VGND VPWR net1429 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[2\]
+ clknet_leaf_61_clk sg13g2_dfrbpq_1
X_6535__187 VPWR VGND net187 sg13g2_tiehi
Xhold270 _1265_ VPWR VGND net1027 sg13g2_dlygate4sd3_1
XFILLER_3_969 VPWR VGND sg13g2_decap_8
XFILLER_49_54 VPWR VGND sg13g2_decap_8
Xhold292 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[3\] VPWR VGND net1049
+ sg13g2_dlygate4sd3_1
Xhold281 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[4\] VPWR VGND net1038
+ sg13g2_dlygate4sd3_1
XFILLER_49_98 VPWR VGND sg13g2_fill_1
XFILLER_19_804 VPWR VGND sg13g2_fill_1
X_6581__141 VPWR VGND net141 sg13g2_tiehi
XFILLER_19_837 VPWR VGND sg13g2_fill_2
XFILLER_34_829 VPWR VGND sg13g2_fill_1
XFILLER_6_741 VPWR VGND sg13g2_decap_8
X_6750__491 VPWR VGND net675 sg13g2_tiehi
XFILLER_2_991 VPWR VGND sg13g2_decap_8
X_4120_ VGND VPWR _1089_ _1088_ _1086_ sg13g2_or2_1
X_4051_ net372 _1041_ _1042_ _1043_ VPWR VGND sg13g2_nor3_1
Xinput5 ui_in[3] net5 VPWR VGND sg13g2_buf_1
XFILLER_36_100 VPWR VGND sg13g2_fill_1
X_6660__62 VPWR VGND net62 sg13g2_tiehi
X_4953_ _1777_ _0617_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[12\]
+ _1783_ VPWR VGND sg13g2_mux2_1
X_3904_ _0630_ _0915_ _0922_ VPWR VGND sg13g2_and2_1
X_4884_ VGND VPWR _1721_ _1723_ _0215_ _1725_ sg13g2_a21oi_1
X_6623_ net99 VGND VPWR _0232_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[8\]
+ clknet_leaf_27_clk sg13g2_dfrbpq_1
X_3835_ _0873_ net552 _0636_ VPWR VGND sg13g2_nand2_1
X_6554_ net168 VGND VPWR net1039 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[4\]
+ clknet_leaf_40_clk sg13g2_dfrbpq_1
X_3766_ _0004_ _0817_ _0818_ _0551_ _0539_ VPWR VGND sg13g2_a22oi_1
X_6485_ net237 VGND VPWR _0094_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].z_sign
+ clknet_leaf_43_clk sg13g2_dfrbpq_2
X_5505_ VGND VPWR _2229_ _2231_ _0328_ _2233_ sg13g2_a21oi_1
X_5436_ _2171_ _2175_ _2176_ VPWR VGND sg13g2_nor2_1
X_3697_ net403 _0685_ net404 _0750_ VPWR VGND sg13g2_nand3_1
X_5367_ VGND VPWR _2109_ _2114_ _2117_ _2112_ sg13g2_a21oi_1
XFILLER_0_906 VPWR VGND sg13g2_decap_8
X_6866__353 VPWR VGND net353 sg13g2_tiehi
X_4318_ _1247_ _1252_ _1246_ _1255_ VPWR VGND sg13g2_nand3_1
X_5298_ _2059_ net415 net1313 VPWR VGND sg13g2_nand2_1
X_4249_ _1196_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[2\]
+ _1195_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_659 VPWR VGND sg13g2_fill_1
XFILLER_24_884 VPWR VGND sg13g2_fill_1
XFILLER_7_527 VPWR VGND sg13g2_fill_1
XFILLER_3_766 VPWR VGND sg13g2_decap_8
XFILLER_46_486 VPWR VGND sg13g2_fill_1
X_3620_ _0673_ _0640_ _0671_ VPWR VGND sg13g2_xnor2_1
X_3551_ VPWR _0621_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[7\] VGND
+ sg13g2_inv_1
X_6270_ net1041 _0605_ _2871_ VPWR VGND net1070 sg13g2_nand3b_1
X_3482_ VPWR _0552_ net889 VGND sg13g2_inv_1
X_5221_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[11\] _1991_ _1996_
+ _1997_ VPWR VGND sg13g2_nor3_1
X_5152_ VGND VPWR _1931_ _1938_ _0269_ _1939_ sg13g2_a21oi_1
X_4103_ _1075_ net532 net834 VPWR VGND sg13g2_xnor2_1
X_5083_ net449 net11 _0257_ VPWR VGND sg13g2_and2_1
X_4034_ _1028_ net551 net885 VPWR VGND sg13g2_nand2b_1
X_6525__197 VPWR VGND net197 sg13g2_tiehi
X_5985_ VGND VPWR net810 _2632_ _0408_ _2633_ sg13g2_a21oi_1
X_4936_ net946 _0544_ _1769_ VPWR VGND sg13g2_nor2_1
X_4867_ _1711_ _0615_ _1710_ VPWR VGND sg13g2_xnor2_1
X_6606_ net116 VGND VPWR _0215_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[4\]
+ clknet_leaf_24_clk sg13g2_dfrbpq_1
X_3818_ _0813_ VPWR _0858_ VGND _0803_ _0805_ sg13g2_o21ai_1
X_4798_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[12\] VPWR _1654_ VGND
+ net536 _1646_ sg13g2_o21ai_1
X_6537_ net185 VGND VPWR net987 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[0\]
+ clknet_leaf_31_clk sg13g2_dfrbpq_1
X_3749_ _0802_ net403 _0801_ VPWR VGND sg13g2_nand2_1
X_6571__151 VPWR VGND net151 sg13g2_tiehi
X_6468_ net259 VGND VPWR net829 u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[7\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_2
X_5419_ _2161_ net1379 _2159_ VPWR VGND sg13g2_xnor2_1
X_6399_ net564 VGND VPWR _0008_ u_angle_cordic_12b_pmod.u_vga_top.clk_div_cnt\[1\]
+ clknet_leaf_65_clk sg13g2_dfrbpq_1
XFILLER_0_703 VPWR VGND sg13g2_decap_8
XFILLER_44_935 VPWR VGND sg13g2_fill_2
XFILLER_12_865 VPWR VGND sg13g2_decap_8
XFILLER_8_825 VPWR VGND sg13g2_decap_8
X_6849__392 VPWR VGND net576 sg13g2_tiehi
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk VPWR VGND sg13g2_buf_8
XFILLER_4_1021 VPWR VGND sg13g2_decap_8
XFILLER_47_795 VPWR VGND sg13g2_fill_1
XFILLER_34_456 VPWR VGND sg13g2_fill_1
XFILLER_21_106 VPWR VGND sg13g2_fill_1
X_5770_ _2456_ net412 net1078 VPWR VGND sg13g2_nand2_1
X_4721_ _1590_ _1583_ _1588_ VPWR VGND sg13g2_nand2_1
X_4652_ _1532_ net1253 net394 VPWR VGND sg13g2_xnor2_1
X_3603_ net403 net408 _0656_ VPWR VGND sg13g2_xor2_1
XFILLER_30_695 VPWR VGND sg13g2_fill_2
Xhold803 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[6\] VPWR VGND net1560
+ sg13g2_dlygate4sd3_1
X_4583_ net1133 net540 _1474_ VPWR VGND sg13g2_xor2_1
X_6322_ net464 net793 _0493_ VPWR VGND sg13g2_and2_1
Xhold814 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[7\] VPWR
+ VGND net1571 sg13g2_dlygate4sd3_1
X_3534_ _0604_ net1525 VPWR VGND sg13g2_inv_2
X_6253_ _2858_ net967 _0543_ VPWR VGND sg13g2_nand2_1
X_3465_ VPWR _0535_ net978 VGND sg13g2_inv_1
X_5204_ VGND VPWR _1976_ _1981_ _0278_ _1982_ sg13g2_a21oi_1
X_6184_ _2802_ net1508 _2804_ VPWR VGND sg13g2_xor2_1
X_5135_ VGND VPWR _1924_ _1923_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[6\]
+ sg13g2_or2_1
X_5066_ _1872_ VPWR _1877_ VGND _1871_ _1873_ sg13g2_o21ai_1
X_4017_ _1014_ _1012_ _1013_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_979 VPWR VGND sg13g2_decap_8
X_5968_ _2625_ _2617_ _2621_ _2624_ VPWR VGND sg13g2_and3_1
X_4919_ net388 VPWR _1755_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[9\]
+ net1173 sg13g2_o21ai_1
X_5899_ _2565_ net1242 _2563_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_68 VPWR VGND sg13g2_fill_1
XFILLER_5_828 VPWR VGND sg13g2_decap_8
X_6393__389 VPWR VGND net573 sg13g2_tiehi
XFILLER_0_522 VPWR VGND sg13g2_fill_1
XFILLER_48_537 VPWR VGND sg13g2_fill_2
XFILLER_17_913 VPWR VGND sg13g2_decap_8
XFILLER_43_275 VPWR VGND sg13g2_fill_2
XFILLER_31_437 VPWR VGND sg13g2_fill_2
X_6679__43 VPWR VGND net43 sg13g2_tiehi
XFILLER_8_699 VPWR VGND sg13g2_fill_1
XFILLER_26_1000 VPWR VGND sg13g2_decap_8
XFILLER_47_570 VPWR VGND sg13g2_fill_1
X_6561__161 VPWR VGND net161 sg13g2_tiehi
X_6871_ net343 VGND VPWR _0480_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[3\]
+ clknet_leaf_11_clk sg13g2_dfrbpq_1
X_5822_ _2497_ _2498_ _2499_ VPWR VGND sg13g2_nor2b_1
X_5753_ _2442_ net517 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[4\]
+ VPWR VGND sg13g2_nand2_1
X_4704_ VGND VPWR _1569_ _1573_ _1575_ net432 sg13g2_a21oi_1
X_5684_ VGND VPWR _2379_ _2383_ _0356_ _2384_ sg13g2_a21oi_1
X_4635_ _1515_ _1516_ _1517_ VPWR VGND sg13g2_nor2b_2
Xhold611 _0316_ VPWR VGND net1368 sg13g2_dlygate4sd3_1
Xhold600 _0097_ VPWR VGND net1357 sg13g2_dlygate4sd3_1
X_4566_ net1038 net539 _1460_ VPWR VGND sg13g2_xor2_1
Xhold622 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[4\]\[2\] VPWR VGND net1379
+ sg13g2_dlygate4sd3_1
XFILLER_2_809 VPWR VGND sg13g2_decap_8
Xhold644 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[7\] VPWR VGND net1401
+ sg13g2_dlygate4sd3_1
Xhold633 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[9\] VPWR VGND net1390
+ sg13g2_dlygate4sd3_1
X_3517_ VPWR _0587_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[11\] VGND
+ sg13g2_inv_1
X_6305_ net462 net764 _0479_ VPWR VGND sg13g2_and2_1
Xhold655 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[6\] VPWR VGND net1412
+ sg13g2_dlygate4sd3_1
Xhold688 _0307_ VPWR VGND net1445 sg13g2_dlygate4sd3_1
Xhold666 _2543_ VPWR VGND net1423 sg13g2_dlygate4sd3_1
Xhold677 _1810_ VPWR VGND net1434 sg13g2_dlygate4sd3_1
X_4497_ _1404_ net1480 _1402_ VPWR VGND sg13g2_xnor2_1
Xhold699 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[3\] VPWR
+ VGND net1456 sg13g2_dlygate4sd3_1
X_6236_ _2845_ net508 net1071 VPWR VGND sg13g2_xnor2_1
X_6167_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[7\] _2788_
+ _2789_ VPWR VGND sg13g2_and2_1
X_5118_ _1907_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[4\]
+ _1909_ VPWR VGND sg13g2_xor2_1
X_6098_ _2730_ net454 _2729_ VPWR VGND sg13g2_nand2_1
X_5049_ net464 VPWR _1863_ VGND _1861_ _1862_ sg13g2_o21ai_1
XFILLER_14_927 VPWR VGND sg13g2_decap_8
XFILLER_25_286 VPWR VGND sg13g2_fill_2
XFILLER_40_245 VPWR VGND sg13g2_fill_2
XFILLER_22_993 VPWR VGND sg13g2_decap_8
XFILLER_49_1000 VPWR VGND sg13g2_decap_8
X_6676__46 VPWR VGND net46 sg13g2_tiehi
XFILLER_1_875 VPWR VGND sg13g2_decap_8
X_6469__257 VPWR VGND net257 sg13g2_tiehi
X_6846__395 VPWR VGND net579 sg13g2_tiehi
XFILLER_48_367 VPWR VGND sg13g2_fill_1
XFILLER_20_919 VPWR VGND sg13g2_decap_8
XFILLER_9_953 VPWR VGND sg13g2_decap_8
XFILLER_13_993 VPWR VGND sg13g2_decap_8
X_4420_ _1339_ net1411 _1337_ VPWR VGND sg13g2_xnor2_1
X_4351_ _1273_ VPWR _1281_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].z_sign
+ _0606_ sg13g2_o21ai_1
X_4282_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[10\] _1224_
+ _1225_ VPWR VGND sg13g2_nor2b_1
Xfanout409 _0641_ net409 VPWR VGND sg13g2_buf_8
X_6021_ net1264 _2661_ _2662_ VPWR VGND sg13g2_and2_1
XFILLER_12_0 VPWR VGND sg13g2_fill_2
X_6923_ net252 VGND VPWR _0518_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[17\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_1
X_6854_ net562 VGND VPWR _0463_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[11\]
+ clknet_leaf_7_clk sg13g2_dfrbpq_2
X_3997_ _0997_ net940 _0995_ VPWR VGND sg13g2_nand2_1
X_6785_ net640 VGND VPWR _0394_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[2\]
+ clknet_leaf_60_clk sg13g2_dfrbpq_1
X_5805_ _2484_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[2\]
+ _2483_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_919 VPWR VGND sg13g2_decap_8
X_5736_ net431 net904 _2429_ _0363_ VPWR VGND sg13g2_nor3_1
X_5667_ net474 VPWR _2370_ VGND _2364_ _2369_ sg13g2_o21ai_1
X_4618_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[2\] _1501_ _1502_
+ VPWR VGND sg13g2_and2_1
X_5598_ net475 VPWR _2311_ VGND _2306_ _2310_ sg13g2_o21ai_1
X_4549_ net760 net436 _0159_ VPWR VGND sg13g2_nor2_1
Xhold463 _1870_ VPWR VGND net1220 sg13g2_dlygate4sd3_1
Xhold441 _0247_ VPWR VGND net1198 sg13g2_dlygate4sd3_1
Xhold452 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[5\] VPWR VGND net1209
+ sg13g2_dlygate4sd3_1
Xhold430 _0233_ VPWR VGND net1187 sg13g2_dlygate4sd3_1
Xhold474 _2275_ VPWR VGND net1231 sg13g2_dlygate4sd3_1
Xhold485 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[0\] VPWR
+ VGND net1242 sg13g2_dlygate4sd3_1
Xhold496 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[6\] VPWR VGND net1253
+ sg13g2_dlygate4sd3_1
X_6219_ _2831_ net508 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[5\]
+ VPWR VGND sg13g2_nand2_1
X_6673__49 VPWR VGND net49 sg13g2_tiehi
XFILLER_38_78 VPWR VGND sg13g2_fill_1
XFILLER_18_518 VPWR VGND sg13g2_fill_2
X_6876__333 VPWR VGND net333 sg13g2_tiehi
XFILLER_14_779 VPWR VGND sg13g2_fill_2
XFILLER_6_923 VPWR VGND sg13g2_decap_8
XFILLER_10_985 VPWR VGND sg13g2_decap_8
X_6551__171 VPWR VGND net171 sg13g2_tiehi
XFILLER_1_672 VPWR VGND sg13g2_decap_8
X_3920_ net450 net776 _0050_ VPWR VGND sg13g2_and2_1
X_3851_ net1019 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[6\] u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[5\]
+ _0883_ VPWR VGND sg13g2_nor3_1
X_3782_ net896 VPWR _0009_ VGND _0826_ _0829_ sg13g2_o21ai_1
X_6570_ net152 VGND VPWR _0179_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[8\]
+ clknet_leaf_26_clk sg13g2_dfrbpq_2
X_5521_ net481 VPWR _2247_ VGND _2243_ _2246_ sg13g2_o21ai_1
X_5452_ _2190_ _0555_ _2188_ VPWR VGND sg13g2_xnor2_1
X_5383_ _2131_ _2130_ _2127_ VPWR VGND sg13g2_nand2b_1
X_4403_ _1322_ net1452 _1324_ VPWR VGND sg13g2_xor2_1
X_4334_ VGND VPWR _1263_ net1027 _0123_ _1267_ sg13g2_a21oi_1
X_6004_ net460 VPWR _2649_ VGND _2647_ _2648_ sg13g2_o21ai_1
X_4265_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[4\] _1202_
+ _1208_ _1210_ VPWR VGND sg13g2_nor3_1
X_4196_ VGND VPWR _0587_ _1137_ _1152_ net534 sg13g2_a21oi_1
X_6906_ net288 VGND VPWR _0501_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[0\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_1
X_6837_ net588 VGND VPWR net1236 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[6\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_10_204 VPWR VGND sg13g2_fill_1
X_6768_ net657 VGND VPWR net1244 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[1\]
+ clknet_leaf_61_clk sg13g2_dfrbpq_1
X_6699_ net740 VGND VPWR _0308_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[8\]
+ clknet_leaf_56_clk sg13g2_dfrbpq_2
X_5719_ _2412_ VPWR _2415_ VGND _2408_ _2413_ sg13g2_o21ai_1
Xhold271 _0123_ VPWR VGND net1028 sg13g2_dlygate4sd3_1
XFILLER_3_948 VPWR VGND sg13g2_decap_8
Xhold260 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[0\] VPWR
+ VGND net1017 sg13g2_dlygate4sd3_1
XFILLER_49_33 VPWR VGND sg13g2_decap_8
Xhold282 _0163_ VPWR VGND net1039 sg13g2_dlygate4sd3_1
Xhold293 _0444_ VPWR VGND net1050 sg13g2_dlygate4sd3_1
X_6843__398 VPWR VGND net582 sg13g2_tiehi
XFILLER_19_849 VPWR VGND sg13g2_fill_2
X_6739__502 VPWR VGND net686 sg13g2_tiehi
XFILLER_41_340 VPWR VGND sg13g2_fill_1
XFILLER_6_720 VPWR VGND sg13g2_decap_8
XFILLER_6_797 VPWR VGND sg13g2_decap_8
XFILLER_2_970 VPWR VGND sg13g2_decap_8
X_4050_ VGND VPWR _1038_ _1039_ _1042_ _1037_ sg13g2_a21oi_1
Xinput6 ui_in[4] net6 VPWR VGND sg13g2_buf_1
XFILLER_25_808 VPWR VGND sg13g2_fill_1
X_4952_ _0226_ net469 _1781_ _1782_ VPWR VGND sg13g2_and3_1
X_4883_ net484 VPWR _1725_ VGND _1721_ _1723_ sg13g2_o21ai_1
X_3903_ _0630_ _0911_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[4\] _0921_ VPWR VGND
+ sg13g2_nand3_1
X_3834_ _0872_ _0539_ net889 VPWR VGND sg13g2_nand2_1
XFILLER_33_885 VPWR VGND sg13g2_fill_1
X_6622_ net100 VGND VPWR net1123 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[7\]
+ clknet_leaf_28_clk sg13g2_dfrbpq_1
X_6553_ net169 VGND VPWR _0162_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[3\]
+ clknet_leaf_39_clk sg13g2_dfrbpq_1
X_3765_ VGND VPWR _0812_ _0816_ _0818_ _0539_ sg13g2_a21oi_1
X_3696_ VGND VPWR _0684_ _0692_ _0749_ _0691_ sg13g2_a21oi_1
X_6484_ net238 VGND VPWR _0093_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[10\]
+ clknet_leaf_43_clk sg13g2_dfrbpq_1
X_5504_ _2233_ net481 _2232_ VPWR VGND sg13g2_nand2_1
X_5435_ _2175_ net1008 _2173_ VPWR VGND sg13g2_xnor2_1
X_5366_ net429 _2115_ _2116_ _0306_ VPWR VGND sg13g2_nor3_1
X_4317_ VGND VPWR net1361 _1253_ _0119_ _1254_ sg13g2_a21oi_1
X_5297_ _2056_ _2057_ _2058_ VPWR VGND sg13g2_nor2_1
X_4248_ _0582_ VPWR _1195_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[0\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[1\] sg13g2_o21ai_1
X_4179_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[10\] _1130_ _1131_
+ _1137_ VPWR VGND sg13g2_nor3_1
X_6541__181 VPWR VGND net181 sg13g2_tiehi
XFILLER_3_745 VPWR VGND sg13g2_decap_8
XFILLER_20_1017 VPWR VGND sg13g2_decap_8
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
XFILLER_18_156 VPWR VGND sg13g2_fill_1
XFILLER_15_885 VPWR VGND sg13g2_decap_8
X_3550_ _0620_ net1546 VPWR VGND sg13g2_inv_2
X_3481_ VPWR _0551_ net929 VGND sg13g2_inv_1
X_5220_ net527 _0571_ _1996_ VPWR VGND sg13g2_nor2_1
X_5151_ net493 VPWR _1939_ VGND _1931_ _1938_ sg13g2_o21ai_1
X_5082_ net449 net10 _0256_ VPWR VGND sg13g2_and2_1
X_4102_ net532 net834 _1074_ VPWR VGND sg13g2_nor2b_1
X_4033_ VGND VPWR _1023_ _1024_ _1027_ _1022_ sg13g2_a21oi_1
XFILLER_37_454 VPWR VGND sg13g2_fill_1
X_5984_ net467 VPWR _2633_ VGND net810 _2632_ sg13g2_o21ai_1
X_4935_ VGND VPWR _1766_ _1767_ _0223_ _1768_ sg13g2_a21oi_1
X_4866_ _0613_ VPWR _1710_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[0\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[1\] sg13g2_o21ai_1
X_6605_ net117 VGND VPWR net1448 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[3\]
+ clknet_leaf_25_clk sg13g2_dfrbpq_1
X_4797_ net536 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[12\] _1646_
+ _1653_ VPWR VGND sg13g2_nor3_1
X_3817_ net553 net866 _0857_ VPWR VGND sg13g2_nor2_1
XFILLER_20_343 VPWR VGND sg13g2_fill_2
X_6536_ net186 VGND VPWR net1288 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[10\]
+ clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_20_376 VPWR VGND sg13g2_fill_1
X_3748_ _0801_ _0753_ _0790_ VPWR VGND sg13g2_nand2_1
X_6467_ net261 VGND VPWR _0076_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[6\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
X_3679_ _0718_ _0638_ _0732_ VPWR VGND sg13g2_xor2_1
X_5418_ _2159_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[4\]\[2\] _2160_
+ VPWR VGND sg13g2_nor2b_1
X_6398_ net565 VGND VPWR _0007_ u_angle_cordic_12b_pmod.u_vga_top.clk_div_cnt\[0\]
+ clknet_leaf_65_clk sg13g2_dfrbpq_1
X_5349_ VGND VPWR _2092_ _2100_ _2102_ net429 sg13g2_a21oi_1
X_6729__512 VPWR VGND net696 sg13g2_tiehi
XFILLER_0_759 VPWR VGND sg13g2_decap_8
XFILLER_46_23 VPWR VGND sg13g2_fill_2
XFILLER_44_947 VPWR VGND sg13g2_fill_2
XFILLER_43_446 VPWR VGND sg13g2_fill_2
X_6736__505 VPWR VGND net689 sg13g2_tiehi
X_6404__372 VPWR VGND net556 sg13g2_tiehi
Xclkbuf_leaf_50_clk clknet_4_11_0_clk clknet_leaf_50_clk VPWR VGND sg13g2_buf_8
XFILLER_8_815 VPWR VGND sg13g2_fill_1
XFILLER_4_1000 VPWR VGND sg13g2_decap_8
XFILLER_22_608 VPWR VGND sg13g2_decap_4
X_4720_ VGND VPWR _1589_ _1588_ _1583_ sg13g2_or2_1
Xclkbuf_leaf_41_clk clknet_4_14_0_clk clknet_leaf_41_clk VPWR VGND sg13g2_buf_8
X_4651_ _1531_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[6\] net393
+ VPWR VGND sg13g2_nand2_1
X_3602_ net408 net403 _0655_ VPWR VGND sg13g2_and2_1
X_4582_ VGND VPWR _1469_ _1471_ _0165_ _1473_ sg13g2_a21oi_1
Xhold804 _0242_ VPWR VGND net1561 sg13g2_dlygate4sd3_1
X_6321_ net463 net784 _0492_ VPWR VGND sg13g2_and2_1
Xhold815 _0383_ VPWR VGND net1572 sg13g2_dlygate4sd3_1
X_3533_ VPWR _0603_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[10\] VGND
+ sg13g2_inv_1
X_6252_ _2857_ net1041 net967 VPWR VGND sg13g2_nand2b_1
X_3464_ VPWR _0534_ net914 VGND sg13g2_inv_1
XFILLER_42_0 VPWR VGND sg13g2_fill_2
X_5203_ net494 VPWR _1982_ VGND _1976_ _1981_ sg13g2_o21ai_1
X_6183_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[9\] _2802_
+ _2803_ VPWR VGND sg13g2_and2_1
X_5134_ VGND VPWR _0566_ _1908_ _1923_ net526 sg13g2_a21oi_1
X_6531__191 VPWR VGND net191 sg13g2_tiehi
XFILLER_29_207 VPWR VGND sg13g2_fill_1
X_5065_ _1876_ net1548 net396 VPWR VGND sg13g2_xnor2_1
X_4016_ _1007_ VPWR _1013_ VGND _1005_ _1006_ sg13g2_o21ai_1
XFILLER_26_936 VPWR VGND sg13g2_fill_1
X_5967_ _2624_ _0581_ _2622_ VPWR VGND sg13g2_xnor2_1
XFILLER_40_405 VPWR VGND sg13g2_fill_1
X_4918_ _1747_ _1749_ _1754_ VPWR VGND sg13g2_nor2b_1
Xclkbuf_leaf_32_clk clknet_4_12_0_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
X_5898_ _2563_ net1242 _2564_ VPWR VGND sg13g2_nor2b_1
XFILLER_32_36 VPWR VGND sg13g2_fill_1
X_4849_ VGND VPWR _1694_ _1695_ _0209_ _1696_ sg13g2_a21oi_1
XFILLER_5_807 VPWR VGND sg13g2_decap_8
XFILLER_10_1027 VPWR VGND sg13g2_fill_2
X_6519_ net203 VGND VPWR net1141 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[7\]
+ clknet_leaf_42_clk sg13g2_dfrbpq_1
XFILLER_28_262 VPWR VGND sg13g2_fill_2
XFILLER_43_232 VPWR VGND sg13g2_fill_2
XFILLER_17_969 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_23_clk clknet_4_7_0_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
Xheichips25_CORDIC_30 VPWR VGND uio_oe[6] sg13g2_tielo
XFILLER_4_895 VPWR VGND sg13g2_decap_8
X_6870_ net345 VGND VPWR _0479_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[2\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_1
X_5821_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[4\] VPWR _2498_
+ VGND _2489_ _2496_ sg13g2_o21ai_1
XFILLER_16_991 VPWR VGND sg13g2_decap_8
X_5752_ VGND VPWR _2437_ _2440_ _0367_ _2441_ sg13g2_a21oi_1
X_6719__522 VPWR VGND net706 sg13g2_tiehi
X_4703_ _1569_ _1573_ _1574_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_14_clk clknet_4_4_0_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
X_5683_ net475 VPWR _2384_ VGND _2379_ _2383_ sg13g2_o21ai_1
X_4634_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[12\] VPWR _1516_ VGND
+ net537 _1514_ sg13g2_o21ai_1
X_4565_ _1459_ _0608_ net1038 VPWR VGND sg13g2_nand2_1
Xhold601 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[4\] VPWR VGND net1358
+ sg13g2_dlygate4sd3_1
Xhold612 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[2\] VPWR
+ VGND net1369 sg13g2_dlygate4sd3_1
Xhold623 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[5\]\[4\] VPWR VGND net1380
+ sg13g2_dlygate4sd3_1
Xhold645 _2317_ VPWR VGND net1402 sg13g2_dlygate4sd3_1
Xhold634 _0309_ VPWR VGND net1391 sg13g2_dlygate4sd3_1
X_3516_ VPWR _0586_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[8\] VGND
+ sg13g2_inv_1
X_6304_ net462 net767 _0478_ VPWR VGND sg13g2_and2_1
Xhold656 _2310_ VPWR VGND net1413 sg13g2_dlygate4sd3_1
Xhold678 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[6\] VPWR
+ VGND net1435 sg13g2_dlygate4sd3_1
Xhold667 _0386_ VPWR VGND net1424 sg13g2_dlygate4sd3_1
X_6392__390 VPWR VGND net574 sg13g2_tiehi
X_4496_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[4\] _1402_
+ _1403_ VPWR VGND sg13g2_nor2_1
Xhold689 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[3\]\[2\] VPWR VGND net1446
+ sg13g2_dlygate4sd3_1
X_6235_ VGND VPWR net417 net1267 _2844_ _2842_ sg13g2_a21oi_1
X_6166_ _2788_ net1371 _2787_ VPWR VGND sg13g2_xnor2_1
X_6726__515 VPWR VGND net699 sg13g2_tiehi
X_6097_ _2727_ VPWR _2729_ VGND _2720_ _2723_ sg13g2_o21ai_1
X_5117_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[4\] _1907_
+ _1908_ VPWR VGND sg13g2_nor2_1
X_5048_ _1862_ net1430 net396 VPWR VGND sg13g2_xnor2_1
XFILLER_27_69 VPWR VGND sg13g2_fill_1
XFILLER_14_906 VPWR VGND sg13g2_decap_8
XFILLER_26_788 VPWR VGND sg13g2_fill_2
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk VPWR VGND sg13g2_buf_8
XFILLER_43_68 VPWR VGND sg13g2_fill_1
XFILLER_22_972 VPWR VGND sg13g2_decap_8
X_6733__508 VPWR VGND net692 sg13g2_tiehi
XFILLER_1_854 VPWR VGND sg13g2_decap_8
XFILLER_29_571 VPWR VGND sg13g2_fill_2
XFILLER_13_972 VPWR VGND sg13g2_decap_8
XFILLER_9_932 VPWR VGND sg13g2_decap_8
X_4350_ _1275_ _1277_ _1280_ VPWR VGND sg13g2_nor2_1
XFILLER_4_692 VPWR VGND sg13g2_decap_8
X_4281_ VGND VPWR _0585_ _1210_ _1224_ net531 sg13g2_a21oi_1
X_6020_ _2661_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[2\]
+ _2660_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_3_clk clknet_4_1_0_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_6922_ net254 VGND VPWR _0517_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[16\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_2
X_6853_ net566 VGND VPWR _0462_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[10\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_2
X_5804_ net413 VPWR _2483_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[0\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[1\] sg13g2_o21ai_1
X_3996_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[0\] _0995_ _0996_
+ VPWR VGND sg13g2_and2_1
X_6784_ net641 VGND VPWR net1250 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[1\]
+ clknet_leaf_61_clk sg13g2_dfrbpq_2
XFILLER_13_38 VPWR VGND sg13g2_fill_1
X_5735_ _2429_ net903 _2425_ _2427_ VPWR VGND sg13g2_and3_1
X_5666_ VPWR _2369_ _2368_ VGND sg13g2_inv_1
X_4617_ _1501_ net1273 _1500_ VPWR VGND sg13g2_xnor2_1
X_5597_ _2310_ net1412 _2308_ VPWR VGND sg13g2_xnor2_1
Xhold420 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[3\] VPWR
+ VGND net1177 sg13g2_dlygate4sd3_1
Xhold453 _2687_ VPWR VGND net1210 sg13g2_dlygate4sd3_1
Xhold442 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[12\] VPWR VGND net1199
+ sg13g2_dlygate4sd3_1
Xhold431 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[1\] VPWR
+ VGND net1188 sg13g2_dlygate4sd3_1
X_4548_ VGND VPWR _1444_ _1445_ _0158_ _1446_ sg13g2_a21oi_1
Xhold464 _0244_ VPWR VGND net1221 sg13g2_dlygate4sd3_1
Xhold486 _2480_ VPWR VGND net1243 sg13g2_dlygate4sd3_1
Xhold475 _0339_ VPWR VGND net1232 sg13g2_dlygate4sd3_1
X_4479_ _1388_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[2\]
+ _1386_ VPWR VGND sg13g2_xnor2_1
X_6218_ VGND VPWR _2826_ _2828_ _0444_ _2830_ sg13g2_a21oi_1
Xhold497 _0177_ VPWR VGND net1254 sg13g2_dlygate4sd3_1
X_6149_ _2773_ _0621_ _2772_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_57 VPWR VGND sg13g2_fill_2
XFILLER_14_758 VPWR VGND sg13g2_fill_2
XFILLER_22_780 VPWR VGND sg13g2_fill_2
XFILLER_6_902 VPWR VGND sg13g2_decap_8
XFILLER_10_964 VPWR VGND sg13g2_decap_8
XFILLER_6_979 VPWR VGND sg13g2_decap_8
XFILLER_1_651 VPWR VGND sg13g2_decap_8
XFILLER_49_622 VPWR VGND sg13g2_fill_1
X_6709__532 VPWR VGND net716 sg13g2_tiehi
XFILLER_0_172 VPWR VGND sg13g2_fill_2
XFILLER_48_121 VPWR VGND sg13g2_fill_2
X_6672__50 VPWR VGND net50 sg13g2_tiehi
XFILLER_36_305 VPWR VGND sg13g2_fill_2
XFILLER_17_585 VPWR VGND sg13g2_decap_4
XFILLER_32_522 VPWR VGND sg13g2_fill_2
X_3850_ _0881_ _0882_ _0024_ VPWR VGND sg13g2_nor2_1
X_3781_ _0828_ net554 _0829_ VPWR VGND _0630_ sg13g2_nand3b_1
X_6716__525 VPWR VGND net709 sg13g2_tiehi
X_5520_ VGND VPWR _2246_ _2245_ _2244_ sg13g2_or2_1
X_5451_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[2\] _2188_
+ _2189_ VPWR VGND sg13g2_and2_1
X_5382_ _0308_ net478 _2129_ _2130_ VPWR VGND sg13g2_and3_1
X_4402_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[3\] _1322_ _1323_
+ VPWR VGND sg13g2_and2_1
X_4333_ _1267_ net502 _1266_ VPWR VGND sg13g2_nand2_1
X_4264_ _1202_ _1208_ _1209_ VPWR VGND sg13g2_nor2_1
X_6003_ _2648_ net514 net1068 VPWR VGND sg13g2_xnor2_1
X_4195_ VGND VPWR _1148_ _1151_ _1149_ _1145_ sg13g2_a21oi_2
X_6905__290 VPWR VGND net290 sg13g2_tiehi
X_6723__518 VPWR VGND net702 sg13g2_tiehi
X_6905_ net290 VGND VPWR net1 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.resetn
+ clknet_leaf_54_clk sg13g2_dfrbpq_2
X_6836_ net589 VGND VPWR net1331 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[5\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_1
X_6767_ net658 VGND VPWR net1016 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[0\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_1
X_5718_ VGND VPWR _2408_ net1450 _0360_ _2414_ sg13g2_a21oi_1
X_3979_ _0980_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[10\] _0947_
+ VPWR VGND sg13g2_xnor2_1
X_6698_ net741 VGND VPWR net1445 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[7\]
+ clknet_leaf_56_clk sg13g2_dfrbpq_1
X_5649_ _2354_ net1240 _2352_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_927 VPWR VGND sg13g2_decap_8
XFILLER_49_12 VPWR VGND sg13g2_decap_8
Xhold250 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[1\] VPWR VGND net1007
+ sg13g2_dlygate4sd3_1
Xhold261 _0185_ VPWR VGND net1018 sg13g2_dlygate4sd3_1
XFILLER_46_1026 VPWR VGND sg13g2_fill_2
Xhold272 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[17\] VPWR VGND net1029
+ sg13g2_dlygate4sd3_1
Xhold283 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[5\] VPWR VGND net1040 sg13g2_dlygate4sd3_1
Xhold294 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[7\] VPWR VGND net1051
+ sg13g2_dlygate4sd3_1
XFILLER_49_89 VPWR VGND sg13g2_decap_8
XFILLER_33_308 VPWR VGND sg13g2_fill_2
XFILLER_41_396 VPWR VGND sg13g2_fill_2
XFILLER_10_794 VPWR VGND sg13g2_fill_2
XFILLER_6_776 VPWR VGND sg13g2_decap_8
X_6414__352 VPWR VGND net352 sg13g2_tiehi
XFILLER_39_6 VPWR VGND sg13g2_fill_2
Xinput7 ui_in[5] net7 VPWR VGND sg13g2_buf_1
XFILLER_18_872 VPWR VGND sg13g2_fill_1
X_4951_ _1782_ _1776_ _1780_ VPWR VGND sg13g2_nand2b_1
XFILLER_17_382 VPWR VGND sg13g2_fill_2
X_3902_ VGND VPWR net901 _0918_ _0920_ net914 sg13g2_a21oi_1
X_4882_ _1721_ _1723_ _1724_ VPWR VGND sg13g2_nor2_1
X_3833_ VGND VPWR net553 _0871_ _0018_ net870 sg13g2_a21oi_1
X_6621_ net101 VGND VPWR _0230_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[6\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_1
X_6552_ net170 VGND VPWR _0161_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[2\]
+ clknet_leaf_39_clk sg13g2_dfrbpq_1
X_3764_ VGND VPWR _0817_ _0816_ _0812_ sg13g2_or2_1
X_3695_ VGND VPWR _0668_ _0695_ _0748_ _0694_ sg13g2_a21oi_1
X_6483_ net239 VGND VPWR net1116 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[9\]
+ clknet_leaf_43_clk sg13g2_dfrbpq_1
X_5503_ VGND VPWR _2232_ _2231_ _2229_ sg13g2_or2_1
X_5434_ _2173_ net1008 _2174_ VPWR VGND sg13g2_nor2b_1
X_5365_ _2109_ _2114_ _2116_ VPWR VGND sg13g2_and2_1
X_4316_ net501 VPWR _1254_ VGND _1252_ _1253_ sg13g2_o21ai_1
X_5296_ _2049_ VPWR _2057_ VGND net528 _0572_ sg13g2_o21ai_1
X_4247_ _1191_ VPWR _1194_ VGND _1187_ _1192_ sg13g2_o21ai_1
X_4178_ _1134_ _1129_ _1133_ _1136_ VPWR VGND sg13g2_a21o_1
X_6819_ net606 VGND VPWR _0428_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[2\]\[1\]
+ clknet_leaf_62_clk sg13g2_dfrbpq_1
XFILLER_13_1014 VPWR VGND sg13g2_decap_8
XFILLER_3_724 VPWR VGND sg13g2_decap_8
X_6706__535 VPWR VGND net719 sg13g2_tiehi
X_6713__528 VPWR VGND net712 sg13g2_tiehi
XFILLER_6_540 VPWR VGND sg13g2_fill_1
X_3480_ VPWR _0550_ net944 VGND sg13g2_inv_1
X_5150_ _1938_ _0568_ _1936_ VPWR VGND sg13g2_xnor2_1
X_4101_ net799 net435 _0084_ VPWR VGND sg13g2_nor2_1
X_5081_ net449 net9 _0255_ VPWR VGND sg13g2_and2_1
X_4032_ _1026_ net885 net376 VPWR VGND sg13g2_nand2_1
XFILLER_37_422 VPWR VGND sg13g2_fill_2
X_5983_ _2632_ net513 net841 VPWR VGND sg13g2_xnor2_1
X_4934_ net483 VPWR _1768_ VGND _1766_ _1767_ sg13g2_o21ai_1
XFILLER_21_812 VPWR VGND sg13g2_fill_1
X_4865_ _1706_ VPWR _1709_ VGND _1702_ _1707_ sg13g2_o21ai_1
X_4796_ _0200_ net483 _1651_ _1652_ VPWR VGND sg13g2_and3_1
X_6604_ net118 VGND VPWR _0213_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[2\]
+ clknet_leaf_26_clk sg13g2_dfrbpq_1
X_3816_ _0016_ _0855_ _0856_ _0550_ _0539_ VPWR VGND sg13g2_a22oi_1
X_3747_ _0792_ VPWR _0800_ VGND _0775_ _0793_ sg13g2_o21ai_1
X_6535_ net187 VGND VPWR net1159 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[3\]
+ clknet_leaf_33_clk sg13g2_dfrbpq_2
X_6466_ net263 VGND VPWR _0075_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[5\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3678_ _0645_ _0703_ _0731_ VPWR VGND sg13g2_nor2_1
X_5417_ _2159_ _0558_ _2158_ VPWR VGND sg13g2_xnor2_1
X_6397_ net567 VGND VPWR net814 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[10\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_1
X_5348_ _2092_ _2100_ _2101_ VPWR VGND sg13g2_nor2_1
XFILLER_0_738 VPWR VGND sg13g2_decap_8
X_5279_ VGND VPWR _2039_ _2041_ _0292_ _2043_ sg13g2_a21oi_1
XFILLER_28_444 VPWR VGND sg13g2_fill_1
XFILLER_8_805 VPWR VGND sg13g2_fill_1
XFILLER_3_543 VPWR VGND sg13g2_fill_2
XFILLER_2_0 VPWR VGND sg13g2_fill_2
Xfanout390 _1722_ net390 VPWR VGND sg13g2_buf_2
XFILLER_19_422 VPWR VGND sg13g2_fill_2
X_4650_ _1528_ _1529_ _1530_ VPWR VGND sg13g2_nor2_1
XFILLER_30_697 VPWR VGND sg13g2_fill_1
X_3601_ _0654_ _0637_ _0653_ VPWR VGND sg13g2_nand2_1
Xinput10 uio_in[0] net10 VPWR VGND sg13g2_buf_1
X_6320_ net464 net779 _0491_ VPWR VGND sg13g2_and2_1
X_4581_ _1473_ net503 _1472_ VPWR VGND sg13g2_nand2_1
Xhold805 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[8\] VPWR VGND net1562
+ sg13g2_dlygate4sd3_1
Xhold816 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[5\] VPWR VGND net1573
+ sg13g2_dlygate4sd3_1
X_3532_ VPWR _0602_ net1441 VGND sg13g2_inv_1
X_6251_ _0451_ net455 _2855_ net1100 VPWR VGND sg13g2_and3_1
X_3463_ VPWR _0533_ net885 VGND sg13g2_inv_1
X_5202_ VPWR _1981_ _1980_ VGND sg13g2_inv_1
X_6182_ _2802_ net1130 _2801_ VPWR VGND sg13g2_xnor2_1
X_5133_ VGND VPWR _1916_ _1921_ _0267_ _1922_ sg13g2_a21oi_1
X_5064_ VGND VPWR _1871_ _1874_ _0245_ _1875_ sg13g2_a21oi_1
X_4015_ net550 net948 _1012_ VPWR VGND sg13g2_xor2_1
X_5966_ _2623_ _0581_ _2622_ VPWR VGND sg13g2_nand2_1
XFILLER_34_970 VPWR VGND sg13g2_fill_2
X_4917_ net388 net1564 _1753_ VPWR VGND sg13g2_xor2_1
X_5897_ _2563_ net1481 _2562_ VPWR VGND sg13g2_xnor2_1
X_4848_ net471 VPWR _1696_ VGND _1694_ _1695_ sg13g2_o21ai_1
X_4779_ _1638_ net1082 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[9\]
+ VPWR VGND sg13g2_xnor2_1
XFILLER_10_1006 VPWR VGND sg13g2_decap_8
X_6518_ net204 VGND VPWR net1193 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[6\]
+ clknet_leaf_40_clk sg13g2_dfrbpq_1
X_6449_ net295 VGND VPWR _0058_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[2\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_2
XFILLER_0_535 VPWR VGND sg13g2_fill_1
XFILLER_44_723 VPWR VGND sg13g2_fill_2
X_6703__538 VPWR VGND net722 sg13g2_tiehi
XFILLER_17_948 VPWR VGND sg13g2_decap_8
XFILLER_29_786 VPWR VGND sg13g2_fill_1
XFILLER_43_277 VPWR VGND sg13g2_fill_1
X_6892__543 VPWR VGND net727 sg13g2_tiehi
XFILLER_31_439 VPWR VGND sg13g2_fill_1
XFILLER_8_613 VPWR VGND sg13g2_fill_2
XFILLER_40_962 VPWR VGND sg13g2_fill_2
XFILLER_22_70 VPWR VGND sg13g2_fill_1
Xheichips25_CORDIC_31 VPWR VGND uio_out[0] sg13g2_tielo
XFILLER_4_874 VPWR VGND sg13g2_decap_8
X_5820_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[4\] _2489_
+ _2496_ _2497_ VPWR VGND sg13g2_nor3_1
XFILLER_16_970 VPWR VGND sg13g2_decap_8
XFILLER_23_929 VPWR VGND sg13g2_decap_8
XFILLER_35_789 VPWR VGND sg13g2_fill_2
X_5751_ net472 VPWR _2441_ VGND _2437_ _2440_ sg13g2_o21ai_1
X_4702_ _1573_ net1438 _1571_ VPWR VGND sg13g2_xnor2_1
X_5682_ _2383_ net1377 _2381_ VPWR VGND sg13g2_xnor2_1
X_4633_ net537 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[12\] _1514_
+ _1515_ VPWR VGND sg13g2_nor3_1
X_4564_ VGND VPWR _1454_ _1457_ _0162_ _1458_ sg13g2_a21oi_1
Xhold602 _0331_ VPWR VGND net1359 sg13g2_dlygate4sd3_1
Xhold624 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[3\] VPWR
+ VGND net1381 sg13g2_dlygate4sd3_1
Xhold635 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[9\] VPWR VGND net1392
+ sg13g2_dlygate4sd3_1
X_3515_ VPWR _0585_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[5\]
+ VGND sg13g2_inv_1
X_6303_ net462 net765 _0477_ VPWR VGND sg13g2_and2_1
Xhold613 _1362_ VPWR VGND net1370 sg13g2_dlygate4sd3_1
Xhold657 _0344_ VPWR VGND net1414 sg13g2_dlygate4sd3_1
Xhold646 _0345_ VPWR VGND net1403 sg13g2_dlygate4sd3_1
Xhold668 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[6\] VPWR
+ VGND net1425 sg13g2_dlygate4sd3_1
Xhold679 _2606_ VPWR VGND net1436 sg13g2_dlygate4sd3_1
X_6234_ _2842_ _2843_ _0447_ VPWR VGND sg13g2_nor2_1
X_4495_ VGND VPWR _0601_ _1387_ _1402_ net543 sg13g2_a21oi_1
X_6165_ net507 _2780_ _2787_ VPWR VGND sg13g2_nor2_1
X_5116_ VGND VPWR _0565_ _1892_ _1907_ net526 sg13g2_a21oi_1
X_6096_ _2720_ _2723_ _2727_ _2728_ VPWR VGND sg13g2_nor3_1
X_5047_ _1861_ _1857_ _1859_ VPWR VGND sg13g2_nand2_1
XFILLER_27_37 VPWR VGND sg13g2_fill_2
X_5949_ _2605_ VPWR _2608_ VGND _2602_ _2606_ sg13g2_o21ai_1
XFILLER_22_951 VPWR VGND sg13g2_decap_8
XFILLER_40_247 VPWR VGND sg13g2_fill_1
XFILLER_21_483 VPWR VGND sg13g2_fill_1
XFILLER_1_833 VPWR VGND sg13g2_decap_8
XFILLER_1_1015 VPWR VGND sg13g2_decap_8
XFILLER_17_756 VPWR VGND sg13g2_fill_1
XFILLER_9_911 VPWR VGND sg13g2_decap_8
XFILLER_13_951 VPWR VGND sg13g2_decap_8
XFILLER_31_258 VPWR VGND sg13g2_fill_1
XFILLER_12_461 VPWR VGND sg13g2_fill_2
X_6517__205 VPWR VGND net205 sg13g2_tiehi
XFILLER_9_988 VPWR VGND sg13g2_decap_8
X_4280_ _1220_ VPWR _1223_ VGND _1217_ _1221_ sg13g2_o21ai_1
X_6921_ net256 VGND VPWR net855 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[15\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_2
X_6852_ net568 VGND VPWR _0461_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[9\]
+ clknet_leaf_7_clk sg13g2_dfrbpq_2
X_6424__332 VPWR VGND net332 sg13g2_tiehi
X_5803_ VGND VPWR _2473_ _2478_ _2482_ net1428 sg13g2_a21oi_1
X_3995_ net550 net924 _0995_ VPWR VGND sg13g2_xor2_1
X_6783_ net642 VGND VPWR net1511 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[0\]
+ clknet_leaf_61_clk sg13g2_dfrbpq_2
X_5734_ VGND VPWR _2425_ _2427_ _2428_ net903 sg13g2_a21oi_1
X_5665_ _2366_ net1230 _2368_ VPWR VGND sg13g2_xor2_1
X_4616_ net538 _1499_ _1500_ VPWR VGND sg13g2_nor2_1
Xhold410 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[4\] VPWR VGND net1167
+ sg13g2_dlygate4sd3_1
X_5596_ _2309_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[6\] _2308_
+ VPWR VGND sg13g2_nand2_1
X_4547_ net498 VPWR _1446_ VGND _1444_ _1445_ sg13g2_o21ai_1
Xhold454 _0419_ VPWR VGND net1211 sg13g2_dlygate4sd3_1
Xhold443 _0120_ VPWR VGND net1200 sg13g2_dlygate4sd3_1
Xhold432 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[7\] VPWR VGND net1189
+ sg13g2_dlygate4sd3_1
Xhold421 _0182_ VPWR VGND net1178 sg13g2_dlygate4sd3_1
Xhold487 _0377_ VPWR VGND net1244 sg13g2_dlygate4sd3_1
Xhold476 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[12\] VPWR VGND net1233
+ sg13g2_dlygate4sd3_1
Xhold465 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[6\] VPWR VGND net1222
+ sg13g2_dlygate4sd3_1
X_4478_ VGND VPWR net411 _1385_ _1387_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[2\]
+ sg13g2_a21oi_1
Xhold498 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[3\] VPWR VGND net1255
+ sg13g2_dlygate4sd3_1
X_6217_ _2830_ net462 _2829_ VPWR VGND sg13g2_nand2_1
X_6148_ VGND VPWR net416 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[6\]
+ _2772_ _2765_ sg13g2_a21oi_1
X_6079_ _2713_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[9\]
+ _2712_ VPWR VGND sg13g2_xnor2_1
XFILLER_41_534 VPWR VGND sg13g2_fill_1
XFILLER_16_1012 VPWR VGND sg13g2_decap_8
XFILLER_10_943 VPWR VGND sg13g2_decap_8
XFILLER_6_958 VPWR VGND sg13g2_decap_8
XFILLER_5_435 VPWR VGND sg13g2_fill_1
XFILLER_23_1027 VPWR VGND sg13g2_fill_2
XFILLER_44_372 VPWR VGND sg13g2_fill_1
X_3780_ net863 net1001 net983 _0827_ _0828_ VPWR VGND sg13g2_nor4_1
XFILLER_13_781 VPWR VGND sg13g2_fill_1
X_5450_ _2188_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[10\] _2187_
+ VPWR VGND sg13g2_xnor2_1
X_4401_ _1322_ _0603_ _1321_ VPWR VGND sg13g2_xnor2_1
X_5381_ _2130_ _2124_ _2128_ VPWR VGND sg13g2_nand2_1
X_4332_ VGND VPWR _1266_ _1265_ _1263_ sg13g2_or2_1
X_4263_ net531 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[3\]
+ _1208_ VPWR VGND sg13g2_nor2b_1
X_6002_ _2645_ VPWR _2647_ VGND net514 _0588_ sg13g2_o21ai_1
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk VPWR VGND sg13g2_buf_8
X_4194_ VGND VPWR _1145_ _1149_ _0100_ _1150_ sg13g2_a21oi_1
X_6904_ net250 VGND VPWR _0521_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[0\].z_sign
+ clknet_leaf_2_clk sg13g2_dfrbpq_2
X_6835_ net590 VGND VPWR net1050 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[4\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_1
X_3978_ _0979_ _0951_ _0978_ VPWR VGND sg13g2_xnor2_1
X_6766_ net659 VGND VPWR net827 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].z_sign
+ clknet_leaf_47_clk sg13g2_dfrbpq_2
X_5717_ net476 VPWR _2414_ VGND _2408_ _2413_ sg13g2_o21ai_1
X_6697_ net742 VGND VPWR _0306_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[6\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_2
X_5648_ _2353_ net1240 _2352_ VPWR VGND sg13g2_nand2_1
X_5579_ net515 _0595_ _2286_ _2294_ VPWR VGND sg13g2_nor3_1
XFILLER_3_906 VPWR VGND sg13g2_decap_8
Xhold262 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[7\] VPWR VGND net1019 sg13g2_dlygate4sd3_1
Xhold251 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[0\] VPWR
+ VGND net1008 sg13g2_dlygate4sd3_1
Xhold240 _0147_ VPWR VGND net997 sg13g2_dlygate4sd3_1
Xhold284 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[0\]\[0\] VPWR VGND net1041
+ sg13g2_dlygate4sd3_1
Xhold273 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[6\] VPWR VGND net1030 sg13g2_dlygate4sd3_1
Xhold295 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].y_shr\[0\] VPWR
+ VGND net1052 sg13g2_dlygate4sd3_1
XFILLER_49_68 VPWR VGND sg13g2_decap_8
XFILLER_18_306 VPWR VGND sg13g2_fill_1
XFILLER_45_103 VPWR VGND sg13g2_fill_2
X_6507__215 VPWR VGND net215 sg13g2_tiehi
XFILLER_42_887 VPWR VGND sg13g2_fill_2
X_6438__309 VPWR VGND net309 sg13g2_tiehi
X_6514__208 VPWR VGND net208 sg13g2_tiehi
XFILLER_6_755 VPWR VGND sg13g2_decap_8
XFILLER_5_265 VPWR VGND sg13g2_fill_1
XFILLER_46_8 VPWR VGND sg13g2_fill_2
XFILLER_49_464 VPWR VGND sg13g2_fill_2
Xinput8 ui_in[6] net8 VPWR VGND sg13g2_buf_1
XFILLER_18_851 VPWR VGND sg13g2_fill_2
XFILLER_45_681 VPWR VGND sg13g2_fill_1
X_4950_ _1781_ _1780_ _1776_ VPWR VGND sg13g2_nand2b_1
XFILLER_17_372 VPWR VGND sg13g2_fill_1
X_4881_ _1723_ net1167 net389 VPWR VGND sg13g2_xnor2_1
X_3901_ VGND VPWR net901 _0918_ _0038_ _0919_ sg13g2_a21oi_1
X_3832_ _0871_ _0865_ _0869_ VPWR VGND sg13g2_xnor2_1
X_6620_ net102 VGND VPWR net1113 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[5\]
+ clknet_leaf_28_clk sg13g2_dfrbpq_1
X_6551_ net171 VGND VPWR _0160_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[1\]
+ clknet_leaf_39_clk sg13g2_dfrbpq_1
X_3763_ _0815_ _0814_ _0816_ VPWR VGND sg13g2_xor2_1
X_5502_ net1074 net524 _2231_ VPWR VGND sg13g2_xor2_1
X_3694_ _0652_ _0746_ _0747_ VPWR VGND sg13g2_and2_1
X_6482_ net240 VGND VPWR net1152 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[8\]
+ clknet_leaf_43_clk sg13g2_dfrbpq_1
X_5433_ _2173_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[8\] _2172_
+ VPWR VGND sg13g2_xnor2_1
X_5364_ _2109_ _2114_ _2115_ VPWR VGND sg13g2_nor2_1
X_4315_ _1234_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[10\] _1251_
+ _1253_ VPWR VGND sg13g2_a21o_1
X_5295_ _2051_ _2053_ _2056_ VPWR VGND sg13g2_nor2_1
X_4246_ VGND VPWR _1187_ _1192_ _0109_ _1193_ sg13g2_a21oi_1
X_4177_ VGND VPWR _1129_ net1364 _0098_ _1135_ sg13g2_a21oi_1
XFILLER_27_125 VPWR VGND sg13g2_fill_1
XFILLER_28_637 VPWR VGND sg13g2_fill_1
X_6838__403 VPWR VGND net587 sg13g2_tiehi
XFILLER_35_26 VPWR VGND sg13g2_fill_1
XFILLER_36_670 VPWR VGND sg13g2_fill_1
X_6818_ net607 VGND VPWR _0427_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[2\]\[0\]
+ clknet_leaf_62_clk sg13g2_dfrbpq_1
X_6749_ net676 VGND VPWR _0358_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[3\]
+ clknet_leaf_56_clk sg13g2_dfrbpq_2
XFILLER_3_703 VPWR VGND sg13g2_decap_8
Xfanout550 net551 net550 VPWR VGND sg13g2_buf_1
X_6627__95 VPWR VGND net95 sg13g2_tiehi
XFILLER_34_629 VPWR VGND sg13g2_fill_1
XFILLER_42_673 VPWR VGND sg13g2_fill_1
XFILLER_30_802 VPWR VGND sg13g2_fill_2
XFILLER_29_1011 VPWR VGND sg13g2_decap_8
X_4100_ net498 net798 _0083_ VPWR VGND sg13g2_and2_1
X_5080_ net448 net8 _0254_ VPWR VGND sg13g2_and2_1
X_4031_ _1021_ VPWR _0062_ VGND net373 _1025_ sg13g2_o21ai_1
X_5982_ net513 net841 _2631_ VPWR VGND sg13g2_nor2b_1
X_4933_ _1767_ net1215 net388 VPWR VGND sg13g2_xnor2_1
XFILLER_33_662 VPWR VGND sg13g2_fill_2
X_4864_ VGND VPWR _1702_ _1707_ _0212_ _1708_ sg13g2_a21oi_1
X_4795_ _1652_ _1644_ _1650_ VPWR VGND sg13g2_nand2_1
X_3815_ net552 _0812_ _0856_ VPWR VGND sg13g2_and2_1
XFILLER_20_345 VPWR VGND sg13g2_fill_1
X_6603_ net119 VGND VPWR net1045 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[1\]
+ clknet_leaf_27_clk sg13g2_dfrbpq_1
X_3746_ _0798_ _0797_ _0799_ VPWR VGND sg13g2_xor2_1
X_6534_ net188 VGND VPWR _0143_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[2\]
+ clknet_leaf_33_clk sg13g2_dfrbpq_2
X_6465_ net265 VGND VPWR _0074_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[4\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_1
X_5416_ net521 _2157_ _2158_ VPWR VGND sg13g2_nor2_1
X_3677_ _0729_ VPWR _0730_ VGND _0727_ _0728_ sg13g2_o21ai_1
X_6396_ net569 VGND VPWR net836 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[9\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
X_5347_ _2098_ _2099_ _2100_ VPWR VGND sg13g2_nor2b_1
XFILLER_0_717 VPWR VGND sg13g2_decap_8
X_5278_ _2043_ net496 _2042_ VPWR VGND sg13g2_nand2_1
XFILLER_47_209 VPWR VGND sg13g2_fill_2
X_4229_ net496 VPWR _1180_ VGND _1178_ _1179_ sg13g2_o21ai_1
X_6504__218 VPWR VGND net218 sg13g2_tiehi
XFILLER_28_478 VPWR VGND sg13g2_fill_2
X_6624__98 VPWR VGND net98 sg13g2_tiehi
XFILLER_12_802 VPWR VGND sg13g2_fill_2
XFILLER_24_640 VPWR VGND sg13g2_fill_2
XFILLER_12_824 VPWR VGND sg13g2_fill_2
XFILLER_12_879 VPWR VGND sg13g2_decap_8
XFILLER_8_839 VPWR VGND sg13g2_decap_8
Xfanout380 _1934_ net380 VPWR VGND sg13g2_buf_8
Xfanout391 net392 net391 VPWR VGND sg13g2_buf_8
Xinput11 uio_in[1] net11 VPWR VGND sg13g2_buf_1
X_3600_ net408 net409 _0653_ VPWR VGND sg13g2_xor2_1
X_4580_ VGND VPWR _1472_ _1471_ _1469_ sg13g2_or2_1
X_3531_ VPWR _0601_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[3\]
+ VGND sg13g2_inv_1
XFILLER_7_883 VPWR VGND sg13g2_decap_8
Xhold817 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[9\] VPWR VGND net1574
+ sg13g2_dlygate4sd3_1
Xhold806 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[5\] VPWR VGND net1563
+ sg13g2_dlygate4sd3_1
X_6250_ net417 VPWR _2856_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[9\]
+ net1099 sg13g2_o21ai_1
X_3462_ VPWR _0532_ net803 VGND sg13g2_inv_1
X_6455__283 VPWR VGND net283 sg13g2_tiehi
X_5201_ _1978_ net1245 _1980_ VPWR VGND sg13g2_xor2_1
X_6828__413 VPWR VGND net597 sg13g2_tiehi
X_6181_ net510 _2795_ _2801_ VPWR VGND sg13g2_nor2_1
X_5132_ net492 VPWR _1922_ VGND _1916_ _1921_ sg13g2_o21ai_1
X_6863__359 VPWR VGND net359 sg13g2_tiehi
XFILLER_28_0 VPWR VGND sg13g2_fill_1
X_5063_ net465 VPWR _1875_ VGND _1871_ _1874_ sg13g2_o21ai_1
XFILLER_38_732 VPWR VGND sg13g2_fill_1
X_4014_ net948 net549 _1011_ VPWR VGND sg13g2_and2_1
XFILLER_25_415 VPWR VGND sg13g2_fill_1
XFILLER_37_264 VPWR VGND sg13g2_fill_1
X_5965_ _2615_ net513 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[12\]
+ _2622_ VPWR VGND sg13g2_mux2_1
X_4916_ _1752_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[10\] net388
+ VPWR VGND sg13g2_nand2_1
X_5896_ net413 VPWR _2562_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[2\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[3\] sg13g2_o21ai_1
X_6835__406 VPWR VGND net590 sg13g2_tiehi
XFILLER_34_993 VPWR VGND sg13g2_fill_2
X_4847_ _1688_ _1693_ _1695_ VPWR VGND sg13g2_and2_1
XFILLER_20_142 VPWR VGND sg13g2_fill_1
XFILLER_20_175 VPWR VGND sg13g2_fill_1
X_4778_ net1082 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[9\] _1637_
+ VPWR VGND sg13g2_nor2b_1
X_3729_ _0782_ _0774_ _0780_ VPWR VGND sg13g2_xnor2_1
X_6517_ net205 VGND VPWR _0126_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[5\]
+ clknet_leaf_40_clk sg13g2_dfrbpq_1
X_6448_ net297 VGND VPWR net925 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[1\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_2
XFILLER_0_503 VPWR VGND sg13g2_fill_2
X_6379_ VGND VPWR _2860_ _2862_ _0455_ net421 sg13g2_a21oi_1
XFILLER_0_514 VPWR VGND sg13g2_fill_2
XFILLER_44_702 VPWR VGND sg13g2_fill_2
XFILLER_16_415 VPWR VGND sg13g2_fill_1
XFILLER_17_927 VPWR VGND sg13g2_decap_8
XFILLER_44_757 VPWR VGND sg13g2_fill_1
XFILLER_19_1010 VPWR VGND sg13g2_decap_8
XFILLER_25_982 VPWR VGND sg13g2_decap_8
XFILLER_11_153 VPWR VGND sg13g2_fill_1
XFILLER_4_853 VPWR VGND sg13g2_decap_8
Xheichips25_CORDIC_32 VPWR VGND uio_out[1] sg13g2_tielo
XFILLER_26_1014 VPWR VGND sg13g2_decap_8
XFILLER_47_562 VPWR VGND sg13g2_fill_2
X_5750_ _2438_ _2439_ _2440_ VPWR VGND sg13g2_nor2b_1
X_4701_ _1571_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[2\] _1572_
+ VPWR VGND sg13g2_nor2b_1
X_5681_ _2382_ net1377 _2381_ VPWR VGND sg13g2_nand2_1
X_4632_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[11\] _1507_ _1514_
+ VPWR VGND sg13g2_nor2b_1
X_4563_ net502 VPWR _1458_ VGND _1454_ _1457_ sg13g2_o21ai_1
Xhold603 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[11\] VPWR VGND net1360
+ sg13g2_dlygate4sd3_1
Xhold625 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[2\] VPWR VGND net1382
+ sg13g2_dlygate4sd3_1
X_6302_ VGND VPWR _2870_ _2887_ _0473_ _2894_ sg13g2_a21oi_1
Xhold636 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[2\] VPWR VGND net1393
+ sg13g2_dlygate4sd3_1
Xhold614 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[9\] VPWR VGND net1371
+ sg13g2_dlygate4sd3_1
X_3514_ VPWR _0584_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[2\]
+ VGND sg13g2_inv_1
X_4494_ _1396_ VPWR _1401_ VGND _1393_ _1397_ sg13g2_o21ai_1
Xhold658 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[4\] VPWR VGND net1415
+ sg13g2_dlygate4sd3_1
Xhold669 _2784_ VPWR VGND net1426 sg13g2_dlygate4sd3_1
Xhold647 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[5\] VPWR VGND net1404
+ sg13g2_dlygate4sd3_1
X_6233_ net455 VPWR _2843_ VGND _2840_ _2841_ sg13g2_o21ai_1
X_6164_ _2784_ _2778_ _2783_ _2786_ VPWR VGND sg13g2_a21o_1
X_5115_ _1902_ VPWR _1906_ VGND _1899_ _1903_ sg13g2_o21ai_1
X_6095_ _2727_ _0624_ _2725_ VPWR VGND sg13g2_xnor2_1
X_5046_ _1860_ _1859_ _0242_ VPWR VGND sg13g2_nor2b_2
X_5948_ VGND VPWR _2602_ net1436 _0397_ _2607_ sg13g2_a21oi_1
XFILLER_22_930 VPWR VGND sg13g2_decap_8
X_5879_ _2547_ net1486 _2549_ VPWR VGND sg13g2_xor2_1
XFILLER_21_451 VPWR VGND sg13g2_fill_2
X_6401__377 VPWR VGND net561 sg13g2_tiehi
XFILLER_49_1014 VPWR VGND sg13g2_decap_8
XFILLER_1_812 VPWR VGND sg13g2_decap_8
XFILLER_1_889 VPWR VGND sg13g2_decap_8
X_6900__551 VPWR VGND net735 sg13g2_tiehi
XFILLER_31_204 VPWR VGND sg13g2_fill_1
X_6818__423 VPWR VGND net607 sg13g2_tiehi
XFILLER_13_930 VPWR VGND sg13g2_decap_8
XFILLER_9_967 VPWR VGND sg13g2_decap_8
X_6825__416 VPWR VGND net600 sg13g2_tiehi
X_6920_ net258 VGND VPWR _0515_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[14\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_1
X_6851_ net570 VGND VPWR _0460_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[8\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_2
XFILLER_23_705 VPWR VGND sg13g2_fill_2
XFILLER_35_543 VPWR VGND sg13g2_fill_2
X_5802_ net1243 _2481_ _0377_ VPWR VGND sg13g2_nor2b_1
X_3994_ _0994_ net924 net549 VPWR VGND sg13g2_nand2_1
X_6782_ net643 VGND VPWR _0391_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[3\]\[2\]
+ clknet_leaf_61_clk sg13g2_dfrbpq_1
X_5733_ VGND VPWR u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[8\]
+ _2416_ _2427_ _2426_ sg13g2_a21oi_1
X_6832__409 VPWR VGND net593 sg13g2_tiehi
X_5664_ _2367_ net1230 _2366_ VPWR VGND sg13g2_nand2_1
XFILLER_30_270 VPWR VGND sg13g2_fill_1
X_4615_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[8\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[9\]
+ _1499_ VPWR VGND sg13g2_nor2_1
X_5595_ _2308_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[6\]
+ _2307_ VPWR VGND sg13g2_xnor2_1
Xhold411 _0216_ VPWR VGND net1168 sg13g2_dlygate4sd3_1
Xhold400 _0333_ VPWR VGND net1157 sg13g2_dlygate4sd3_1
X_4546_ _1445_ net1262 net385 VPWR VGND sg13g2_xnor2_1
Xhold422 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.up VPWR VGND net1179 sg13g2_dlygate4sd3_1
Xhold444 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[2\] VPWR
+ VGND net1201 sg13g2_dlygate4sd3_1
Xhold433 _1537_ VPWR VGND net1190 sg13g2_dlygate4sd3_1
Xhold477 _0312_ VPWR VGND net1234 sg13g2_dlygate4sd3_1
Xhold466 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[2\] VPWR VGND net1223
+ sg13g2_dlygate4sd3_1
X_4477_ _1386_ net411 _1385_ VPWR VGND sg13g2_nand2_1
Xhold455 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[4\] VPWR VGND net1212
+ sg13g2_dlygate4sd3_1
Xhold499 _2090_ VPWR VGND net1256 sg13g2_dlygate4sd3_1
Xhold488 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[5\]\[3\] VPWR VGND net1245
+ sg13g2_dlygate4sd3_1
X_6216_ VGND VPWR _2829_ _2828_ _2826_ sg13g2_or2_1
X_6147_ VPWR _2771_ _2770_ VGND sg13g2_inv_1
X_6681__41 VPWR VGND net41 sg13g2_tiehi
XFILLER_38_59 VPWR VGND sg13g2_fill_1
X_6078_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[8\] net416
+ _2706_ _2712_ VPWR VGND sg13g2_a21o_1
X_5029_ _1847_ _1845_ _1841_ VPWR VGND sg13g2_nand2b_1
XFILLER_10_922 VPWR VGND sg13g2_decap_8
XFILLER_6_937 VPWR VGND sg13g2_decap_8
XFILLER_10_999 VPWR VGND sg13g2_decap_8
XFILLER_5_469 VPWR VGND sg13g2_fill_2
XFILLER_1_686 VPWR VGND sg13g2_decap_8
XFILLER_48_123 VPWR VGND sg13g2_fill_1
XFILLER_0_174 VPWR VGND sg13g2_fill_1
XFILLER_23_1006 VPWR VGND sg13g2_decap_8
XFILLER_36_307 VPWR VGND sg13g2_fill_1
XFILLER_9_786 VPWR VGND sg13g2_fill_2
X_4400_ net410 VPWR _1321_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[9\]
+ _1312_ sg13g2_o21ai_1
X_5380_ VGND VPWR _2129_ _2128_ _2124_ sg13g2_or2_1
X_4331_ _1265_ net542 net1026 VPWR VGND sg13g2_xnor2_1
XFILLER_5_63 VPWR VGND sg13g2_fill_2
X_4262_ _1204_ VPWR _1207_ VGND _1201_ _1205_ sg13g2_o21ai_1
X_6001_ VGND VPWR _2643_ _2644_ _0411_ _2646_ sg13g2_a21oi_1
X_4193_ net495 VPWR _1150_ VGND _1145_ _1149_ sg13g2_o21ai_1
XFILLER_28_808 VPWR VGND sg13g2_fill_1
XFILLER_39_167 VPWR VGND sg13g2_fill_1
X_6903_ net738 VGND VPWR _0520_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[10\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
X_6834_ net591 VGND VPWR _0443_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[3\]
+ clknet_leaf_11_clk sg13g2_dfrbpq_1
XFILLER_35_395 VPWR VGND sg13g2_fill_1
X_6765_ net660 VGND VPWR net1129 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[10\]
+ clknet_leaf_47_clk sg13g2_dfrbpq_1
X_3977_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[11\] _0948_ _0978_
+ VPWR VGND sg13g2_nor2b_1
X_5716_ _2413_ net1449 _2411_ VPWR VGND sg13g2_xnor2_1
X_6696_ net743 VGND VPWR net1418 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[5\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_2
X_5647_ _2352_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[4\] _2351_
+ VPWR VGND sg13g2_xnor2_1
X_5578_ VGND VPWR _2284_ _2291_ _2293_ _2289_ sg13g2_a21oi_1
X_4529_ net384 net1477 _1428_ _1431_ VPWR VGND sg13g2_a21o_1
Xhold252 _0301_ VPWR VGND net1009 sg13g2_dlygate4sd3_1
XFILLER_2_406 VPWR VGND sg13g2_fill_1
Xhold230 _0146_ VPWR VGND net987 sg13g2_dlygate4sd3_1
Xhold241 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[0\] VPWR VGND net998
+ sg13g2_dlygate4sd3_1
XFILLER_46_1028 VPWR VGND sg13g2_fill_1
Xhold296 _0237_ VPWR VGND net1053 sg13g2_dlygate4sd3_1
Xhold285 _0469_ VPWR VGND net1042 sg13g2_dlygate4sd3_1
Xhold263 _0891_ VPWR VGND net1020 sg13g2_dlygate4sd3_1
Xhold274 _0889_ VPWR VGND net1031 sg13g2_dlygate4sd3_1
XFILLER_49_47 VPWR VGND sg13g2_decap_8
X_6808__433 VPWR VGND net617 sg13g2_tiehi
X_6815__426 VPWR VGND net610 sg13g2_tiehi
XFILLER_6_701 VPWR VGND sg13g2_decap_4
XFILLER_6_734 VPWR VGND sg13g2_decap_8
XFILLER_10_796 VPWR VGND sg13g2_fill_1
XFILLER_2_984 VPWR VGND sg13g2_decap_8
XFILLER_49_421 VPWR VGND sg13g2_fill_2
X_6822__419 VPWR VGND net603 sg13g2_tiehi
Xinput9 ui_in[7] net9 VPWR VGND sg13g2_buf_1
X_4880_ _1716_ net536 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[10\]
+ _1722_ VPWR VGND sg13g2_mux2_1
X_3900_ net443 VPWR _0919_ VGND net901 _0918_ sg13g2_o21ai_1
XFILLER_32_332 VPWR VGND sg13g2_fill_1
X_3831_ _0869_ _0865_ _0870_ VPWR VGND sg13g2_nor2b_1
X_6550_ net172 VGND VPWR _0159_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[0\]
+ clknet_leaf_38_clk sg13g2_dfrbpq_1
X_3762_ VGND VPWR _0807_ _0810_ _0815_ _0805_ sg13g2_a21oi_1
X_5501_ _2230_ net418 net1074 VPWR VGND sg13g2_nand2_1
X_3693_ _0744_ _0698_ _0746_ VPWR VGND sg13g2_xor2_1
X_6481_ net241 VGND VPWR net1176 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[7\]
+ clknet_leaf_43_clk sg13g2_dfrbpq_1
X_5432_ VGND VPWR net418 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[7\]
+ _2172_ _2165_ sg13g2_a21oi_1
X_5363_ VPWR _2114_ _2113_ VGND sg13g2_inv_1
X_4314_ _1252_ net1360 _1233_ VPWR VGND sg13g2_xnor2_1
X_5294_ net435 _2054_ _2055_ _0295_ VPWR VGND sg13g2_nor3_1
X_4245_ net479 VPWR _1193_ VGND _1187_ _1192_ sg13g2_o21ai_1
X_4176_ net495 VPWR _1135_ VGND _1129_ _1134_ sg13g2_o21ai_1
Xclkbuf_leaf_62_clk clknet_4_2_0_clk clknet_leaf_62_clk VPWR VGND sg13g2_buf_8
X_6817_ net608 VGND VPWR net1132 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[12\]
+ clknet_leaf_9_clk sg13g2_dfrbpq_2
XFILLER_23_343 VPWR VGND sg13g2_fill_2
X_6873__339 VPWR VGND net339 sg13g2_tiehi
X_6748_ net677 VGND VPWR _0357_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[2\]
+ clknet_leaf_55_clk sg13g2_dfrbpq_1
X_6679_ net43 VGND VPWR _0288_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[0\]
+ clknet_leaf_37_clk sg13g2_dfrbpq_1
X_6437__310 VPWR VGND net310 sg13g2_tiehi
XFILLER_3_759 VPWR VGND sg13g2_decap_8
Xfanout540 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].z_sign net540
+ VPWR VGND sg13g2_buf_8
Xfanout551 net1179 net551 VPWR VGND sg13g2_buf_1
X_6444__303 VPWR VGND net303 sg13g2_tiehi
Xclkbuf_leaf_53_clk clknet_4_10_0_clk clknet_leaf_53_clk VPWR VGND sg13g2_buf_8
X_6520__202 VPWR VGND net202 sg13g2_tiehi
XFILLER_42_696 VPWR VGND sg13g2_fill_2
XFILLER_15_899 VPWR VGND sg13g2_decap_8
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk VPWR VGND sg13g2_buf_8
XFILLER_2_781 VPWR VGND sg13g2_decap_8
X_4030_ _1025_ _1023_ _1024_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_424 VPWR VGND sg13g2_fill_1
XFILLER_18_671 VPWR VGND sg13g2_fill_2
X_5981_ net810 net427 _0407_ VPWR VGND sg13g2_nor2_1
X_4932_ _1766_ _1755_ _1764_ _1765_ VPWR VGND sg13g2_and3_1
XFILLER_24_129 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_44_clk clknet_4_14_0_clk clknet_leaf_44_clk VPWR VGND sg13g2_buf_8
XFILLER_36_1027 VPWR VGND sg13g2_fill_2
X_4863_ net483 VPWR _1708_ VGND _1702_ _1707_ sg13g2_o21ai_1
X_6602_ net120 VGND VPWR net1000 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[0\]
+ clknet_leaf_27_clk sg13g2_dfrbpq_1
X_4794_ VGND VPWR _1651_ _1650_ _1644_ sg13g2_or2_1
X_3814_ _0788_ _0799_ _0811_ _0855_ VPWR VGND sg13g2_or3_1
XFILLER_21_858 VPWR VGND sg13g2_fill_1
X_3745_ _0785_ VPWR _0798_ VGND _0772_ _0786_ sg13g2_o21ai_1
X_6533_ net189 VGND VPWR _0142_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[1\]
+ clknet_leaf_32_clk sg13g2_dfrbpq_2
X_6464_ net267 VGND VPWR _0073_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[3\]
+ clknet_leaf_11_clk sg13g2_dfrbpq_2
X_5415_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[4\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[5\]
+ _2157_ VPWR VGND sg13g2_nor2_1
X_3676_ _0637_ VPWR _0729_ VGND _0638_ _0639_ sg13g2_o21ai_1
X_6395_ net571 VGND VPWR net930 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[5\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
X_5346_ VGND VPWR _2099_ _2097_ net1505 sg13g2_or2_1
X_5277_ VGND VPWR _2042_ _2041_ _2039_ sg13g2_or2_1
X_4228_ VGND VPWR net1300 net382 _1179_ _1177_ sg13g2_a21oi_1
X_6805__436 VPWR VGND net620 sg13g2_tiehi
X_4159_ _1120_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[6\]\[1\] _1118_
+ VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_35_clk clknet_4_12_0_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
XFILLER_23_140 VPWR VGND sg13g2_fill_1
XFILLER_24_696 VPWR VGND sg13g2_fill_2
X_6812__429 VPWR VGND net613 sg13g2_tiehi
XFILLER_11_62 VPWR VGND sg13g2_fill_2
XFILLER_11_84 VPWR VGND sg13g2_fill_1
XFILLER_4_1014 VPWR VGND sg13g2_decap_8
Xfanout381 _1233_ net381 VPWR VGND sg13g2_buf_8
Xfanout392 _1660_ net392 VPWR VGND sg13g2_buf_8
XFILLER_19_424 VPWR VGND sg13g2_fill_1
XFILLER_46_276 VPWR VGND sg13g2_fill_1
XFILLER_35_939 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_26_clk clknet_4_13_0_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
Xinput12 uio_in[2] net12 VPWR VGND sg13g2_buf_1
XFILLER_30_688 VPWR VGND sg13g2_fill_2
XFILLER_11_891 VPWR VGND sg13g2_decap_8
X_3530_ VPWR _0600_ net541 VGND sg13g2_inv_1
Xhold807 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[10\] VPWR VGND net1564
+ sg13g2_dlygate4sd3_1
XFILLER_7_862 VPWR VGND sg13g2_decap_8
Xhold818 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[8\] VPWR VGND net1575
+ sg13g2_dlygate4sd3_1
X_3461_ VPWR _0531_ net856 VGND sg13g2_inv_1
X_5200_ _1979_ net1245 _1978_ VPWR VGND sg13g2_nand2_1
X_6180_ _2798_ _2793_ _2797_ _2800_ VPWR VGND sg13g2_a21o_2
X_5131_ VPWR _1921_ _1920_ VGND sg13g2_inv_1
X_5062_ _1874_ net1260 net395 VPWR VGND sg13g2_xnor2_1
X_4013_ _1010_ net948 net376 VPWR VGND sg13g2_nand2_1
XFILLER_38_700 VPWR VGND sg13g2_fill_2
X_5964_ net425 _2619_ _2620_ _0399_ VPWR VGND sg13g2_nor3_1
Xclkbuf_leaf_17_clk clknet_4_4_0_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
X_4915_ VGND VPWR _1749_ _1750_ _0220_ _1751_ sg13g2_a21oi_1
X_5895_ _2558_ VPWR _2561_ VGND _2554_ _2559_ sg13g2_o21ai_1
X_4846_ _1694_ net1201 net392 VPWR VGND sg13g2_xnor2_1
X_4777_ VPWR VGND _0613_ net436 _1636_ net1142 _0197_ _1632_ sg13g2_a221oi_1
X_6516_ net206 VGND VPWR net1081 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[4\]
+ clknet_leaf_40_clk sg13g2_dfrbpq_1
X_3728_ _0774_ _0780_ _0781_ VPWR VGND sg13g2_nor2b_1
X_6434__313 VPWR VGND net313 sg13g2_tiehi
X_6447_ net299 VGND VPWR _0056_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[0\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_2
X_3659_ _0712_ _0709_ _0710_ VPWR VGND sg13g2_xnor2_1
X_6378_ net878 net442 _0521_ VPWR VGND sg13g2_and2_1
X_5329_ _2078_ _2083_ _2084_ VPWR VGND sg13g2_nor2b_1
X_6510__212 VPWR VGND net212 sg13g2_tiehi
XFILLER_48_519 VPWR VGND sg13g2_fill_1
XFILLER_44_714 VPWR VGND sg13g2_fill_1
XFILLER_16_405 VPWR VGND sg13g2_fill_1
XFILLER_17_906 VPWR VGND sg13g2_decap_8
X_6441__306 VPWR VGND net306 sg13g2_tiehi
XFILLER_25_961 VPWR VGND sg13g2_decap_8
X_6619__103 VPWR VGND net103 sg13g2_tiehi
XFILLER_11_143 VPWR VGND sg13g2_fill_1
XFILLER_12_666 VPWR VGND sg13g2_fill_2
XFILLER_4_832 VPWR VGND sg13g2_decap_8
Xheichips25_CORDIC_33 VPWR VGND uio_out[2] sg13g2_tielo
XFILLER_19_298 VPWR VGND sg13g2_fill_1
X_5680_ _2381_ net1334 _2380_ VPWR VGND sg13g2_xnor2_1
X_4700_ _1571_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[2\]
+ _1570_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_452 VPWR VGND sg13g2_fill_1
X_4631_ VGND VPWR u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[3\] _1509_
+ _1513_ _1512_ sg13g2_a21oi_1
X_4562_ _1455_ _1456_ _1457_ VPWR VGND sg13g2_nor2b_1
Xhold626 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[3\] VPWR VGND net1383
+ sg13g2_dlygate4sd3_1
X_6301_ _2894_ net444 _2871_ VPWR VGND sg13g2_nand2_1
Xhold615 _2722_ VPWR VGND net1372 sg13g2_dlygate4sd3_1
X_3513_ VPWR _0583_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[1\] VGND
+ sg13g2_inv_1
Xhold604 _1252_ VPWR VGND net1361 sg13g2_dlygate4sd3_1
X_4493_ _1396_ _1398_ _1400_ VPWR VGND sg13g2_and2_1
Xhold659 _0343_ VPWR VGND net1416 sg13g2_dlygate4sd3_1
Xhold637 _1897_ VPWR VGND net1394 sg13g2_dlygate4sd3_1
Xclkbuf_leaf_6_clk clknet_4_4_0_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
X_6232_ _2840_ _2841_ _2842_ VPWR VGND sg13g2_and2_1
Xhold648 _0113_ VPWR VGND net1405 sg13g2_dlygate4sd3_1
XFILLER_40_0 VPWR VGND sg13g2_fill_2
X_6163_ VGND VPWR _2778_ net1426 _0434_ _2785_ sg13g2_a21oi_1
X_6094_ _2726_ net1130 _2725_ VPWR VGND sg13g2_nand2_1
X_5114_ _1904_ _1905_ _0265_ VPWR VGND sg13g2_nor2b_1
X_6841__400 VPWR VGND net584 sg13g2_tiehi
X_5045_ net470 VPWR _1860_ VGND _1856_ _1858_ sg13g2_o21ai_1
X_6802__439 VPWR VGND net623 sg13g2_tiehi
XFILLER_27_39 VPWR VGND sg13g2_fill_1
X_5947_ net459 VPWR _2607_ VGND _2602_ _2606_ sg13g2_o21ai_1
X_5878_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[11\] _2547_ _2548_
+ VPWR VGND sg13g2_and2_1
XFILLER_22_986 VPWR VGND sg13g2_decap_8
X_4829_ _1678_ _1679_ _1668_ _1680_ VPWR VGND sg13g2_nand3_1
XFILLER_1_868 VPWR VGND sg13g2_decap_8
X_6922__254 VPWR VGND net254 sg13g2_tiehi
XFILLER_13_986 VPWR VGND sg13g2_decap_8
XFILLER_9_946 VPWR VGND sg13g2_decap_8
Xhold1 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[9\] VPWR VGND net758
+ sg13g2_dlygate4sd3_1
X_6850_ net575 VGND VPWR _0459_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[7\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_2
X_5801_ VGND VPWR _2473_ _2479_ _2481_ net424 sg13g2_a21oi_1
X_6781_ net644 VGND VPWR net1148 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[3\]\[1\]
+ clknet_leaf_61_clk sg13g2_dfrbpq_1
X_5732_ VGND VPWR u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[7\]
+ _2415_ _2426_ _2416_ sg13g2_a21oi_1
X_6500__222 VPWR VGND net222 sg13g2_tiehi
X_3993_ _0993_ net924 net376 VPWR VGND sg13g2_nand2_1
X_5663_ _2366_ net1412 _2365_ VPWR VGND sg13g2_xnor2_1
X_4614_ _1495_ VPWR _1498_ VGND _1491_ _1496_ sg13g2_o21ai_1
X_5594_ net412 VPWR _2307_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[5\]
+ _2295_ sg13g2_o21ai_1
Xhold401 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[3\] VPWR
+ VGND net1158 sg13g2_dlygate4sd3_1
X_4545_ _1444_ _1434_ _1442_ _1443_ VPWR VGND sg13g2_and3_1
Xhold423 _0055_ VPWR VGND net1180 sg13g2_dlygate4sd3_1
Xhold445 _1698_ VPWR VGND net1202 sg13g2_dlygate4sd3_1
Xhold434 _0178_ VPWR VGND net1191 sg13g2_dlygate4sd3_1
Xhold412 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[10\] VPWR VGND net1169
+ sg13g2_dlygate4sd3_1
Xhold478 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[6\] VPWR VGND net1235
+ sg13g2_dlygate4sd3_1
X_4476_ VGND VPWR _1385_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[1\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[0\] sg13g2_or2_1
Xhold456 _0175_ VPWR VGND net1213 sg13g2_dlygate4sd3_1
Xhold467 _1390_ VPWR VGND net1224 sg13g2_dlygate4sd3_1
Xhold489 _0278_ VPWR VGND net1246 sg13g2_dlygate4sd3_1
X_6215_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[4\] net508 _2828_
+ VPWR VGND sg13g2_xor2_1
X_6146_ _2767_ VPWR _2770_ VGND _2764_ _2768_ sg13g2_o21ai_1
X_6609__113 VPWR VGND net113 sg13g2_tiehi
X_6077_ _0422_ net453 net1320 _2711_ VPWR VGND sg13g2_and3_1
X_5028_ _1846_ _1841_ _1845_ VPWR VGND sg13g2_nand2b_1
XFILLER_10_901 VPWR VGND sg13g2_decap_8
X_6616__106 VPWR VGND net106 sg13g2_tiehi
XFILLER_6_916 VPWR VGND sg13g2_decap_8
XFILLER_10_978 VPWR VGND sg13g2_decap_8
X_6883__319 VPWR VGND net319 sg13g2_tiehi
XFILLER_0_131 VPWR VGND sg13g2_fill_2
XFILLER_1_665 VPWR VGND sg13g2_decap_8
XFILLER_32_569 VPWR VGND sg13g2_fill_1
XFILLER_9_743 VPWR VGND sg13g2_fill_2
XFILLER_12_282 VPWR VGND sg13g2_fill_1
X_6831__410 VPWR VGND net594 sg13g2_tiehi
X_4330_ _1264_ net542 net1026 VPWR VGND sg13g2_nand2_1
XFILLER_5_982 VPWR VGND sg13g2_decap_8
X_4261_ VGND VPWR _1201_ _1205_ _0111_ _1206_ sg13g2_a21oi_1
X_6000_ _2646_ net460 _2645_ VPWR VGND sg13g2_nand2_1
X_4192_ _1147_ net1398 _1149_ VPWR VGND sg13g2_xor2_1
X_6902_ net737 VGND VPWR _0530_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[9\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
X_6833_ net592 VGND VPWR _0442_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[2\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_1
X_6764_ net661 VGND VPWR _0373_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[9\]
+ clknet_leaf_30_clk sg13g2_dfrbpq_1
X_3976_ _0954_ _0975_ _0950_ _0977_ VPWR VGND _0976_ sg13g2_nand4_1
X_6695_ net744 VGND VPWR _0304_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[4\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_1
X_5715_ _2412_ net1449 _2411_ VPWR VGND sg13g2_nand2_1
X_5646_ net515 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[3\] _2351_
+ VPWR VGND sg13g2_nor2b_1
Xhold220 _1492_ VPWR VGND net977 sg13g2_dlygate4sd3_1
X_5577_ VGND VPWR _2284_ _2291_ _0341_ _2292_ sg13g2_a21oi_1
X_4528_ net385 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[9\] _1430_
+ VPWR VGND sg13g2_xor2_1
Xhold253 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[3\]\[0\] VPWR VGND net1010
+ sg13g2_dlygate4sd3_1
Xhold242 _1703_ VPWR VGND net999 sg13g2_dlygate4sd3_1
Xhold231 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[0\] VPWR VGND net988
+ sg13g2_dlygate4sd3_1
XFILLER_49_26 VPWR VGND sg13g2_decap_8
Xhold286 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[0\].y_shr\[10\] VPWR
+ VGND net1043 sg13g2_dlygate4sd3_1
Xhold264 _0027_ VPWR VGND net1021 sg13g2_dlygate4sd3_1
Xhold275 _0026_ VPWR VGND net1032 sg13g2_dlygate4sd3_1
X_4459_ _1365_ _1368_ _1371_ VPWR VGND sg13g2_nor2_1
Xhold297 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[4\]\[0\] VPWR VGND net1054
+ sg13g2_dlygate4sd3_1
X_6639__83 VPWR VGND net83 sg13g2_tiehi
X_6129_ net452 VPWR _2756_ VGND _2751_ _2755_ sg13g2_o21ai_1
XFILLER_10_720 VPWR VGND sg13g2_fill_2
XFILLER_5_201 VPWR VGND sg13g2_fill_2
XFILLER_30_50 VPWR VGND sg13g2_fill_1
XFILLER_30_61 VPWR VGND sg13g2_fill_1
XFILLER_2_963 VPWR VGND sg13g2_decap_8
XFILLER_7_1023 VPWR VGND sg13g2_decap_4
XFILLER_49_466 VPWR VGND sg13g2_fill_1
XFILLER_36_138 VPWR VGND sg13g2_fill_2
X_3830_ _0869_ _0862_ _0863_ _0687_ _0636_ VPWR VGND sg13g2_a22oi_1
X_3761_ _0814_ _0802_ _0813_ VPWR VGND sg13g2_xnor2_1
XFILLER_13_591 VPWR VGND sg13g2_fill_1
X_5500_ VGND VPWR net852 _2227_ _2229_ _2226_ sg13g2_a21oi_1
X_3692_ _0698_ _0715_ _0743_ _0745_ VPWR VGND sg13g2_nor3_1
X_6480_ net242 VGND VPWR _0089_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[6\]
+ clknet_leaf_42_clk sg13g2_dfrbpq_1
X_5431_ _2167_ VPWR _2171_ VGND _2164_ _2169_ sg13g2_o21ai_1
X_5362_ _2113_ net1541 _2111_ VPWR VGND sg13g2_xnor2_1
X_4313_ net437 net1528 _1251_ _0118_ VPWR VGND sg13g2_nor3_1
X_5293_ _2055_ _2049_ _2051_ _2053_ VPWR VGND sg13g2_and3_1
X_4244_ _1192_ _0583_ _1190_ VPWR VGND sg13g2_xnor2_1
X_4175_ _1132_ net1363 _1134_ VPWR VGND sg13g2_xor2_1
X_6606__116 VPWR VGND net116 sg13g2_tiehi
X_6636__86 VPWR VGND net86 sg13g2_tiehi
X_6816_ net609 VGND VPWR _0425_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[11\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_2
X_6747_ net678 VGND VPWR net1378 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[1\]
+ clknet_leaf_55_clk sg13g2_dfrbpq_2
X_3959_ _0960_ _0958_ _0959_ VPWR VGND sg13g2_nand2_1
XFILLER_13_1028 VPWR VGND sg13g2_fill_1
X_6678_ net44 VGND VPWR net1316 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[10\]
+ clknet_leaf_50_clk sg13g2_dfrbpq_2
X_6613__109 VPWR VGND net109 sg13g2_tiehi
X_5629_ _2338_ net1467 _2336_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_738 VPWR VGND sg13g2_decap_8
Xfanout530 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].z_sign net530
+ VPWR VGND sg13g2_buf_8
Xfanout541 net542 net541 VPWR VGND sg13g2_buf_8
Xfanout552 u_angle_cordic_12b_pmod.u_vga_top.pixel_clk_en net552 VPWR VGND sg13g2_buf_8
X_6821__420 VPWR VGND net604 sg13g2_tiehi
XFILLER_42_631 VPWR VGND sg13g2_fill_1
XFILLER_42_620 VPWR VGND sg13g2_fill_2
XFILLER_15_845 VPWR VGND sg13g2_fill_1
XFILLER_41_93 VPWR VGND sg13g2_fill_2
XFILLER_2_760 VPWR VGND sg13g2_decap_8
XFILLER_1_281 VPWR VGND sg13g2_fill_1
X_6633__89 VPWR VGND net89 sg13g2_tiehi
X_5980_ net467 net773 _0406_ VPWR VGND sg13g2_and2_1
X_4931_ net388 VPWR _1765_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[10\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[11\] sg13g2_o21ai_1
XFILLER_18_683 VPWR VGND sg13g2_fill_1
XFILLER_36_1017 VPWR VGND sg13g2_fill_1
X_4862_ _1707_ _0614_ _1705_ VPWR VGND sg13g2_xnor2_1
X_6601_ net121 VGND VPWR net1203 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].y_shr\[10\]
+ clknet_leaf_25_clk sg13g2_dfrbpq_2
X_3813_ VGND VPWR net552 _0854_ _0015_ net910 sg13g2_a21oi_1
X_4793_ _1650_ net1470 _1648_ VPWR VGND sg13g2_xnor2_1
X_3744_ _0795_ _0796_ _0797_ VPWR VGND sg13g2_nor2b_1
X_6532_ net190 VGND VPWR _0141_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[0\]
+ clknet_leaf_32_clk sg13g2_dfrbpq_2
X_6463_ net269 VGND VPWR _0072_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[2\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_1
X_3675_ _0718_ VPWR _0728_ VGND _0648_ _0724_ sg13g2_o21ai_1
X_5414_ _2153_ VPWR _2156_ VGND _2149_ _2154_ sg13g2_o21ai_1
X_6394_ net572 VGND VPWR net823 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[0\]\[0\]
+ clknet_leaf_63_clk sg13g2_dfrbpq_2
X_5345_ net1505 _2097_ _2098_ VPWR VGND sg13g2_and2_1
X_5276_ _2041_ net528 net1095 VPWR VGND sg13g2_xnor2_1
X_4227_ _1178_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[5\]
+ net383 VPWR VGND sg13g2_xnor2_1
X_4158_ _1119_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[6\]\[1\] _1118_
+ VPWR VGND sg13g2_nand2_1
X_4089_ VGND VPWR net828 _1066_ _0077_ _1067_ sg13g2_a21oi_1
X_6411__358 VPWR VGND net358 sg13g2_tiehi
Xfanout382 net383 net382 VPWR VGND sg13g2_buf_8
Xfanout393 net394 net393 VPWR VGND sg13g2_buf_8
XFILLER_19_447 VPWR VGND sg13g2_fill_1
XFILLER_28_992 VPWR VGND sg13g2_decap_8
Xinput13 uio_in[3] net13 VPWR VGND sg13g2_buf_1
XFILLER_11_870 VPWR VGND sg13g2_decap_8
XFILLER_7_841 VPWR VGND sg13g2_decap_8
Xhold808 _1757_ VPWR VGND net1565 sg13g2_dlygate4sd3_1
Xhold819 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[3\] VPWR
+ VGND net1576 sg13g2_dlygate4sd3_1
X_5130_ _1920_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[5\] _1918_
+ VPWR VGND sg13g2_xnor2_1
X_5061_ net1260 net395 _1873_ VPWR VGND sg13g2_nor2_1
X_4012_ _1004_ VPWR _0059_ VGND net372 _1009_ sg13g2_o21ai_1
X_6603__119 VPWR VGND net119 sg13g2_tiehi
X_5963_ _2613_ _2611_ _2618_ _2621_ VPWR VGND sg13g2_a21o_1
X_4914_ net484 VPWR _1751_ VGND _1749_ _1750_ sg13g2_o21ai_1
X_5894_ VGND VPWR _2554_ net1147 _0390_ _2560_ sg13g2_a21oi_1
XFILLER_34_995 VPWR VGND sg13g2_fill_1
X_4845_ _0208_ net471 _1692_ _1693_ VPWR VGND sg13g2_and3_1
X_4776_ _1634_ _1635_ _1633_ _1636_ VPWR VGND sg13g2_nand3_1
X_6515_ net207 VGND VPWR _0124_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[3\]
+ clknet_leaf_40_clk sg13g2_dfrbpq_1
X_3727_ _0779_ _0776_ _0780_ VPWR VGND sg13g2_xor2_1
X_6811__430 VPWR VGND net614 sg13g2_tiehi
X_6446_ net301 VGND VPWR net1180 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.up
+ clknet_leaf_17_clk sg13g2_dfrbpq_1
X_3658_ _0709_ _0710_ _0711_ VPWR VGND sg13g2_nor2b_1
X_6377_ VPWR _0518_ _2927_ VGND sg13g2_inv_1
X_3589_ net546 u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[7\] u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[7\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[7\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp\[0\]
+ net544 _0642_ VPWR VGND sg13g2_mux4_1
X_5328_ _2083_ _2082_ _2081_ VPWR VGND sg13g2_nand2b_1
X_5259_ VGND VPWR _2022_ _2027_ _2030_ _2028_ sg13g2_a21oi_1
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk VPWR VGND sg13g2_buf_8
XFILLER_44_704 VPWR VGND sg13g2_fill_1
XFILLER_28_277 VPWR VGND sg13g2_fill_2
X_6890__292 VPWR VGND net292 sg13g2_tiehi
XFILLER_4_811 VPWR VGND sg13g2_decap_8
Xheichips25_CORDIC_34 VPWR VGND uio_out[3] sg13g2_tielo
XFILLER_4_888 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_fill_1
X_6862__361 VPWR VGND net361 sg13g2_tiehi
XFILLER_47_564 VPWR VGND sg13g2_fill_1
XFILLER_47_597 VPWR VGND sg13g2_fill_2
XFILLER_16_984 VPWR VGND sg13g2_decap_8
X_4630_ net433 net1352 _1512_ _0174_ VPWR VGND sg13g2_nor3_1
X_4561_ _1456_ net539 net1419 VPWR VGND sg13g2_nand2b_1
X_6300_ VGND VPWR _2892_ _2893_ _0472_ _2890_ sg13g2_a21oi_1
X_4492_ VGND VPWR _1393_ _1397_ _0149_ _1399_ sg13g2_a21oi_1
Xhold627 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[3\] VPWR VGND net1384
+ sg13g2_dlygate4sd3_1
Xhold616 _0424_ VPWR VGND net1373 sg13g2_dlygate4sd3_1
X_3512_ net531 _0582_ VPWR VGND sg13g2_inv_4
Xhold605 _0119_ VPWR VGND net1362 sg13g2_dlygate4sd3_1
Xhold649 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[4\] VPWR
+ VGND net1406 sg13g2_dlygate4sd3_1
Xhold638 _0264_ VPWR VGND net1395 sg13g2_dlygate4sd3_1
X_6231_ _2837_ VPWR _2841_ VGND _2835_ _2836_ sg13g2_o21ai_1
X_6162_ net453 VPWR _2785_ VGND _2778_ _2784_ sg13g2_o21ai_1
X_5113_ VGND VPWR _1899_ _1903_ _1905_ net430 sg13g2_a21oi_1
X_6093_ _2724_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[11\]
+ _2725_ VPWR VGND sg13g2_xor2_1
X_5044_ _1859_ _1856_ _1858_ VPWR VGND sg13g2_nand2_1
XFILLER_38_575 VPWR VGND sg13g2_fill_2
X_5946_ _2606_ net1435 _2604_ VPWR VGND sg13g2_xnor2_1
X_5877_ _2546_ VPWR _2547_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[10\]
+ _2540_ sg13g2_o21ai_1
XFILLER_22_965 VPWR VGND sg13g2_decap_8
X_4828_ net391 VPWR _1679_ VGND net1091 net1515 sg13g2_o21ai_1
X_4759_ net400 net1273 _1620_ _1621_ VPWR VGND sg13g2_a21o_1
X_7478_ hsync_sig net23 VPWR VGND sg13g2_buf_1
X_6429_ net322 VGND VPWR net902 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[7\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_2
XFILLER_0_302 VPWR VGND sg13g2_fill_1
XFILLER_1_847 VPWR VGND sg13g2_decap_8
XFILLER_29_531 VPWR VGND sg13g2_fill_2
XFILLER_9_925 VPWR VGND sg13g2_decap_8
XFILLER_13_965 VPWR VGND sg13g2_decap_8
XFILLER_4_685 VPWR VGND sg13g2_decap_8
Xhold2 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[1\] VPWR VGND net759
+ sg13g2_dlygate4sd3_1
X_6801__440 VPWR VGND net624 sg13g2_tiehi
XFILLER_35_545 VPWR VGND sg13g2_fill_1
X_3992_ _0990_ VPWR _0056_ VGND net940 net372 sg13g2_o21ai_1
X_6780_ net645 VGND VPWR _0389_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[3\]\[0\]
+ clknet_leaf_61_clk sg13g2_dfrbpq_1
X_5800_ _2473_ _2479_ _2480_ VPWR VGND sg13g2_nor2_1
XFILLER_23_707 VPWR VGND sg13g2_fill_1
X_5731_ VGND VPWR _2425_ _2422_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[8\]
+ sg13g2_or2_1
XFILLER_31_762 VPWR VGND sg13g2_fill_2
X_5662_ VGND VPWR _0596_ _2357_ _2365_ net515 sg13g2_a21oi_1
X_4613_ VGND VPWR _1491_ _1496_ _0172_ _1497_ sg13g2_a21oi_1
X_5593_ VGND VPWR _2300_ _2304_ _2306_ _2303_ sg13g2_a21oi_1
Xhold402 _0144_ VPWR VGND net1159 sg13g2_dlygate4sd3_1
X_4544_ net385 VPWR _1443_ VGND net1169 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[11\]
+ sg13g2_o21ai_1
Xhold413 _0157_ VPWR VGND net1170 sg13g2_dlygate4sd3_1
Xhold424 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[3\] VPWR
+ VGND net1181 sg13g2_dlygate4sd3_1
Xhold435 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[6\] VPWR VGND net1192
+ sg13g2_dlygate4sd3_1
Xhold446 _0210_ VPWR VGND net1203 sg13g2_dlygate4sd3_1
X_6214_ _2827_ net417 net1329 VPWR VGND sg13g2_nand2_1
Xhold468 _1391_ VPWR VGND net1225 sg13g2_dlygate4sd3_1
X_4475_ _1381_ VPWR _1384_ VGND _1377_ _1382_ sg13g2_o21ai_1
Xhold457 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[6\] VPWR VGND net1214
+ sg13g2_dlygate4sd3_1
Xhold479 _0446_ VPWR VGND net1236 sg13g2_dlygate4sd3_1
X_6145_ VGND VPWR _2764_ _2768_ _0432_ _2769_ sg13g2_a21oi_1
X_6076_ _2704_ _2700_ _2709_ _2711_ VPWR VGND sg13g2_a21o_1
X_5027_ _1845_ net1500 net396 VPWR VGND sg13g2_xnor2_1
X_5929_ _2591_ net1575 _2590_ VPWR VGND sg13g2_xnor2_1
XFILLER_16_1026 VPWR VGND sg13g2_fill_2
XFILLER_10_957 VPWR VGND sg13g2_decap_8
XFILLER_29_361 VPWR VGND sg13g2_fill_2
XFILLER_17_589 VPWR VGND sg13g2_fill_1
XFILLER_8_221 VPWR VGND sg13g2_fill_1
XFILLER_8_287 VPWR VGND sg13g2_fill_1
XFILLER_9_788 VPWR VGND sg13g2_fill_1
XFILLER_5_961 VPWR VGND sg13g2_decap_8
X_4260_ net479 VPWR _1206_ VGND _1201_ _1205_ sg13g2_o21ai_1
X_4191_ net1398 _1147_ _1148_ VPWR VGND sg13g2_and2_1
X_6901_ net736 VGND VPWR _0529_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[8\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_36_843 VPWR VGND sg13g2_fill_1
X_6832_ net593 VGND VPWR _0441_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[1\]
+ clknet_leaf_28_clk sg13g2_dfrbpq_1
XFILLER_23_548 VPWR VGND sg13g2_fill_1
X_6763_ net662 VGND VPWR _0372_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[8\]
+ clknet_leaf_30_clk sg13g2_dfrbpq_1
X_3975_ _0976_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[12\] _0967_
+ VPWR VGND sg13g2_xnor2_1
X_6694_ net745 VGND VPWR net1257 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[3\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_5714_ _2411_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[12\] _2409_
+ VPWR VGND sg13g2_xnor2_1
X_5645_ net431 net1011 _0351_ VPWR VGND sg13g2_nor2_1
Xhold210 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[0\].y_shr\[0\] VPWR
+ VGND net967 sg13g2_dlygate4sd3_1
X_5576_ net474 VPWR _2292_ VGND _2284_ _2291_ sg13g2_o21ai_1
X_6912__276 VPWR VGND net276 sg13g2_tiehi
X_4527_ _1428_ _1429_ _0154_ VPWR VGND sg13g2_nor2_1
Xhold221 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[3\] VPWR VGND net978 sg13g2_dlygate4sd3_1
Xhold232 _1826_ VPWR VGND net989 sg13g2_dlygate4sd3_1
Xhold243 _0211_ VPWR VGND net1000 sg13g2_dlygate4sd3_1
Xhold287 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[0\] VPWR
+ VGND net1044 sg13g2_dlygate4sd3_1
Xhold276 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[0\] VPWR VGND net1033
+ sg13g2_dlygate4sd3_1
Xhold254 _2350_ VPWR VGND net1011 sg13g2_dlygate4sd3_1
Xhold265 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[14\] VPWR VGND net1022
+ sg13g2_dlygate4sd3_1
X_4458_ VGND VPWR _1368_ _1369_ _0144_ _1370_ sg13g2_a21oi_1
Xhold298 _2150_ VPWR VGND net1055 sg13g2_dlygate4sd3_1
X_6128_ _2755_ net1298 _2753_ VPWR VGND sg13g2_xnor2_1
X_4389_ _1308_ VPWR _1311_ VGND _1304_ _1309_ sg13g2_o21ai_1
X_6059_ net424 _2695_ _2696_ VPWR VGND sg13g2_nor2_1
X_6622__100 VPWR VGND net100 sg13g2_tiehi
XFILLER_14_526 VPWR VGND sg13g2_fill_2
XFILLER_6_769 VPWR VGND sg13g2_decap_8
XFILLER_2_942 VPWR VGND sg13g2_decap_8
XFILLER_49_423 VPWR VGND sg13g2_fill_1
XFILLER_7_1002 VPWR VGND sg13g2_decap_8
XFILLER_39_71 VPWR VGND sg13g2_fill_2
XFILLER_45_662 VPWR VGND sg13g2_fill_1
XFILLER_33_802 VPWR VGND sg13g2_fill_1
X_6421__338 VPWR VGND net338 sg13g2_tiehi
X_3760_ net404 _0636_ _0813_ VPWR VGND sg13g2_xor2_1
X_5430_ VGND VPWR _2164_ _2169_ _0316_ _2170_ sg13g2_a21oi_1
X_3691_ _0715_ _0743_ _0744_ VPWR VGND sg13g2_nor2_1
X_5361_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[6\] _2111_ _2112_
+ VPWR VGND sg13g2_and2_1
X_5292_ VGND VPWR _2049_ _2051_ _2054_ _2053_ sg13g2_a21oi_1
X_4312_ _1246_ _1249_ _1251_ VPWR VGND sg13g2_and2_1
X_4243_ VGND VPWR _1191_ _1190_ _0583_ sg13g2_or2_1
X_4174_ net1363 _1132_ _1133_ VPWR VGND sg13g2_and2_1
X_6465__265 VPWR VGND net265 sg13g2_tiehi
X_6815_ net610 VGND VPWR net1373 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[10\]
+ clknet_leaf_7_clk sg13g2_dfrbpq_2
XFILLER_24_868 VPWR VGND sg13g2_fill_1
X_6746_ net679 VGND VPWR _0355_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[0\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_2
XFILLER_13_1007 VPWR VGND sg13g2_decap_8
X_3958_ _0959_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[5\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt_sum\[5\]
+ VPWR VGND sg13g2_xnor2_1
X_3889_ _0909_ _0910_ _0911_ _0912_ VPWR VGND sg13g2_nor3_1
X_6677_ net45 VGND VPWR net1229 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[5\]
+ clknet_leaf_48_clk sg13g2_dfrbpq_1
X_5628_ _2336_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[10\] _2337_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_3_717 VPWR VGND sg13g2_decap_8
X_5559_ net1231 _2276_ _0339_ VPWR VGND sg13g2_nor2b_1
Xfanout520 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].z_sign net520
+ VPWR VGND sg13g2_buf_8
Xfanout531 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].z_sign net531
+ VPWR VGND sg13g2_buf_8
Xfanout542 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].z_sign net542
+ VPWR VGND sg13g2_buf_8
Xfanout553 net554 net553 VPWR VGND sg13g2_buf_8
XFILLER_26_172 VPWR VGND sg13g2_fill_2
XFILLER_25_40 VPWR VGND sg13g2_fill_1
XFILLER_41_131 VPWR VGND sg13g2_fill_1
XFILLER_42_698 VPWR VGND sg13g2_fill_1
XFILLER_6_500 VPWR VGND sg13g2_fill_2
XFILLER_29_1025 VPWR VGND sg13g2_decap_4
XFILLER_1_260 VPWR VGND sg13g2_fill_2
XFILLER_46_971 VPWR VGND sg13g2_fill_1
X_4930_ _1754_ _1760_ _1753_ _1764_ VPWR VGND sg13g2_nand3_1
X_4861_ VGND VPWR _1706_ _1705_ _0614_ sg13g2_or2_1
X_3812_ _0854_ _0788_ _0799_ VPWR VGND sg13g2_xnor2_1
X_6872__341 VPWR VGND net341 sg13g2_tiehi
X_6600_ net122 VGND VPWR _0209_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].y_shr\[1\]
+ clknet_leaf_26_clk sg13g2_dfrbpq_2
X_4792_ _1649_ net1470 _1648_ VPWR VGND sg13g2_nand2b_1
X_3743_ _0794_ VPWR _0796_ VGND _0781_ _0783_ sg13g2_o21ai_1
X_6531_ net191 VGND VPWR _0140_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[7\]
+ clknet_leaf_31_clk sg13g2_dfrbpq_1
X_6462_ net271 VGND VPWR _0071_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[1\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_2
X_3674_ _0640_ _0726_ _0727_ VPWR VGND sg13g2_nor2b_1
X_6612__110 VPWR VGND net110 sg13g2_tiehi
X_5413_ VGND VPWR _2149_ _2154_ _0314_ _2155_ sg13g2_a21oi_1
X_6393_ net573 VGND VPWR net861 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[0\].y_shr\[0\]
+ clknet_leaf_65_clk sg13g2_dfrbpq_2
X_5344_ _2094_ _2096_ _2097_ VPWR VGND sg13g2_nor2b_1
X_5275_ _2040_ net528 net1095 VPWR VGND sg13g2_nand2_1
X_4226_ net433 _1176_ _1177_ _0105_ VPWR VGND sg13g2_nor3_1
X_4157_ _1118_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[7\] _1117_
+ VPWR VGND sg13g2_xnor2_1
X_4088_ net445 VPWR _1067_ VGND net828 _1066_ sg13g2_o21ai_1
X_6632__90 VPWR VGND net90 sg13g2_tiehi
XFILLER_24_698 VPWR VGND sg13g2_fill_1
X_6729_ net696 VGND VPWR net935 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[0\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_1
XFILLER_11_64 VPWR VGND sg13g2_fill_1
XFILLER_3_558 VPWR VGND sg13g2_fill_2
Xfanout383 _1159_ net383 VPWR VGND sg13g2_buf_8
Xfanout372 net373 net372 VPWR VGND sg13g2_buf_8
Xfanout394 _1522_ net394 VPWR VGND sg13g2_buf_8
XFILLER_14_142 VPWR VGND sg13g2_fill_2
Xinput14 uio_in[4] net14 VPWR VGND sg13g2_buf_1
XFILLER_7_820 VPWR VGND sg13g2_decap_8
Xhold809 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[2\] VPWR
+ VGND net1566 sg13g2_dlygate4sd3_1
XFILLER_7_897 VPWR VGND sg13g2_decap_8
X_5060_ _1872_ net1260 net395 VPWR VGND sg13g2_nand2_1
X_4011_ _1009_ _1005_ _1008_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_702 VPWR VGND sg13g2_fill_1
XFILLER_26_908 VPWR VGND sg13g2_fill_1
X_5962_ VGND VPWR _2611_ _2613_ _2620_ _2618_ sg13g2_a21oi_1
XFILLER_19_982 VPWR VGND sg13g2_decap_8
X_4913_ _1750_ _1745_ _1747_ VPWR VGND sg13g2_nand2_1
X_5893_ net457 VPWR _2560_ VGND _2554_ _2559_ sg13g2_o21ai_1
XFILLER_34_985 VPWR VGND sg13g2_fill_2
X_4844_ _1691_ _1690_ _1689_ _1693_ VPWR VGND sg13g2_a21o_1
X_4775_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[7\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[6\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[5\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[4\]
+ _1635_ VPWR VGND sg13g2_nor4_1
X_6514_ net208 VGND VPWR net1028 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[2\]
+ clknet_leaf_38_clk sg13g2_dfrbpq_1
X_3726_ _0779_ _0777_ _0778_ VPWR VGND sg13g2_nand2_1
X_6445_ net302 VGND VPWR _0054_ u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[11\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_1
X_3657_ _0710_ _0663_ _0665_ VPWR VGND sg13g2_xnor2_1
X_6376_ _2926_ VPWR _2927_ VGND net1029 _2925_ sg13g2_o21ai_1
X_3588_ net546 u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[6\] u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[6\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[6\] net535 net544 _0641_
+ VPWR VGND sg13g2_mux4_1
X_5327_ _2082_ _0556_ _2080_ VPWR VGND sg13g2_nand2_1
X_5258_ _2029_ _2022_ _2027_ _2028_ VPWR VGND sg13g2_and3_1
X_5189_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[5\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[6\]
+ _1969_ VPWR VGND sg13g2_nor2_1
X_4209_ net433 _1162_ _1163_ _0102_ VPWR VGND sg13g2_nor3_1
XFILLER_19_1024 VPWR VGND sg13g2_decap_4
XFILLER_25_996 VPWR VGND sg13g2_decap_8
XFILLER_12_668 VPWR VGND sg13g2_fill_1
Xheichips25_CORDIC_35 VPWR VGND uio_out[4] sg13g2_tielo
Xheichips25_CORDIC_24 VPWR VGND uio_oe[0] sg13g2_tielo
XFILLER_4_867 VPWR VGND sg13g2_decap_8
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
XFILLER_19_278 VPWR VGND sg13g2_fill_1
X_6602__120 VPWR VGND net120 sg13g2_tiehi
XFILLER_34_237 VPWR VGND sg13g2_fill_1
XFILLER_16_963 VPWR VGND sg13g2_decap_8
XFILLER_30_410 VPWR VGND sg13g2_fill_2
X_4560_ net539 net1419 _1455_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_54 VPWR VGND sg13g2_fill_1
Xhold606 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[6\]\[3\] VPWR VGND net1363
+ sg13g2_dlygate4sd3_1
X_3511_ VPWR _0581_ net1531 VGND sg13g2_inv_1
Xhold617 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[4\] VPWR VGND net1374
+ sg13g2_dlygate4sd3_1
X_4491_ _1399_ net486 _1398_ VPWR VGND sg13g2_nand2_1
Xhold639 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[5\] VPWR VGND net1396
+ sg13g2_dlygate4sd3_1
Xhold628 _2290_ VPWR VGND net1385 sg13g2_dlygate4sd3_1
X_6230_ _2840_ net509 net1267 VPWR VGND sg13g2_xnor2_1
X_6161_ _2784_ net1425 _2781_ VPWR VGND sg13g2_xnor2_1
X_5112_ _1899_ _1903_ _1904_ VPWR VGND sg13g2_nor2_1
X_6092_ _2718_ VPWR _2724_ VGND net510 _0625_ sg13g2_o21ai_1
X_5043_ _1858_ net1560 net396 VPWR VGND sg13g2_xnor2_1
XFILLER_25_204 VPWR VGND sg13g2_fill_1
XFILLER_25_215 VPWR VGND sg13g2_fill_2
X_5945_ _2605_ net1435 _2604_ VPWR VGND sg13g2_nand2_1
X_5876_ _2546_ net513 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[10\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_22_944 VPWR VGND sg13g2_decap_8
X_4827_ _1664_ _1665_ _1677_ _1678_ VPWR VGND sg13g2_or3_1
X_4758_ net433 _1619_ _1620_ _0194_ VPWR VGND sg13g2_nor3_1
X_7477_ u_angle_cordic_12b_pmod.u_vga_top.vsync net20 VPWR VGND sg13g2_buf_1
X_3709_ _0762_ _0761_ _0681_ VPWR VGND sg13g2_nand2b_1
X_4689_ _1562_ net993 net1017 VPWR VGND sg13g2_nand2_1
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
X_6428_ net324 VGND VPWR net943 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[6\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_2
XFILLER_1_826 VPWR VGND sg13g2_decap_8
X_6359_ net975 _2913_ _2916_ VPWR VGND sg13g2_nor2_1
XFILLER_29_510 VPWR VGND sg13g2_fill_1
XFILLER_1_1008 VPWR VGND sg13g2_decap_8
XFILLER_29_587 VPWR VGND sg13g2_fill_2
XFILLER_13_944 VPWR VGND sg13g2_decap_8
XFILLER_9_904 VPWR VGND sg13g2_decap_8
X_6452__289 VPWR VGND net289 sg13g2_tiehi
Xhold3 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[0\] VPWR VGND net760
+ sg13g2_dlygate4sd3_1
XFILLER_0_892 VPWR VGND sg13g2_decap_8
X_3991_ _0992_ net372 VPWR VGND sg13g2_inv_2
X_5730_ VGND VPWR _2422_ net1118 _0362_ _2424_ sg13g2_a21oi_1
XFILLER_43_590 VPWR VGND sg13g2_fill_1
X_5661_ VGND VPWR _2356_ _2361_ _2364_ _2360_ sg13g2_a21oi_1
X_4612_ net498 VPWR _1497_ VGND _1491_ _1496_ sg13g2_o21ai_1
X_5592_ VGND VPWR _2300_ _2304_ _0343_ _2305_ sg13g2_a21oi_1
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk VPWR VGND sg13g2_buf_8
X_4543_ _1433_ _1435_ _1439_ _1442_ VPWR VGND sg13g2_or3_1
Xhold403 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[1\] VPWR VGND net1160
+ sg13g2_dlygate4sd3_1
Xhold425 _0284_ VPWR VGND net1182 sg13g2_dlygate4sd3_1
Xhold414 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[9\] VPWR VGND net1171
+ sg13g2_dlygate4sd3_1
Xhold436 _0127_ VPWR VGND net1193 sg13g2_dlygate4sd3_1
Xhold458 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[12\] VPWR VGND net1215
+ sg13g2_dlygate4sd3_1
X_6431__318 VPWR VGND net318 sg13g2_tiehi
X_6213_ VGND VPWR net508 net1049 _2826_ _2825_ sg13g2_a21oi_1
Xhold447 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[4\] VPWR VGND net1204
+ sg13g2_dlygate4sd3_1
X_4474_ VGND VPWR _1377_ _1382_ _0147_ _1383_ sg13g2_a21oi_1
Xhold469 _0148_ VPWR VGND net1226 sg13g2_dlygate4sd3_1
X_6144_ net453 VPWR _2769_ VGND _2764_ _2768_ sg13g2_o21ai_1
XFILLER_38_18 VPWR VGND sg13g2_fill_2
X_6075_ _2704_ _2709_ net1319 _2710_ VPWR VGND sg13g2_nand3_1
X_5026_ _1844_ net1500 net395 VPWR VGND sg13g2_nand2_1
X_5928_ VGND VPWR net413 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[7\]
+ _2590_ _2583_ sg13g2_a21oi_1
XFILLER_16_1005 VPWR VGND sg13g2_decap_8
XFILLER_10_936 VPWR VGND sg13g2_decap_8
X_5859_ _2532_ _2525_ _2530_ VPWR VGND sg13g2_nand2b_1
XFILLER_0_133 VPWR VGND sg13g2_fill_1
XFILLER_29_340 VPWR VGND sg13g2_fill_2
XFILLER_45_877 VPWR VGND sg13g2_fill_1
XFILLER_9_745 VPWR VGND sg13g2_fill_1
XFILLER_5_940 VPWR VGND sg13g2_decap_8
X_4190_ _1147_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[11\] _1146_
+ VPWR VGND sg13g2_xnor2_1
X_6648__74 VPWR VGND net74 sg13g2_tiehi
X_6900_ net735 VGND VPWR _0528_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[7\]
+ clknet_leaf_6_clk sg13g2_dfrbpq_1
X_6831_ net594 VGND VPWR net762 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[0\]
+ clknet_leaf_28_clk sg13g2_dfrbpq_1
XFILLER_23_527 VPWR VGND sg13g2_fill_2
XFILLER_23_538 VPWR VGND sg13g2_fill_1
X_6762_ net663 VGND VPWR net1079 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[7\]
+ clknet_leaf_30_clk sg13g2_dfrbpq_1
X_3974_ _0969_ _0972_ _0973_ _0974_ _0975_ VPWR VGND sg13g2_nor4_1
X_6693_ net746 VGND VPWR net1518 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[2\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_5713_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[12\] _2409_ _2410_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_31_571 VPWR VGND sg13g2_fill_2
X_5644_ _2350_ net1010 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[3\]
+ VPWR VGND sg13g2_xnor2_1
Xhold211 _2858_ VPWR VGND net968 sg13g2_dlygate4sd3_1
X_5575_ VPWR _2291_ net1385 VGND sg13g2_inv_1
Xhold200 _2911_ VPWR VGND net957 sg13g2_dlygate4sd3_1
X_4526_ net498 VPWR _1429_ VGND _1425_ _1427_ sg13g2_o21ai_1
Xhold244 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[9\] VPWR VGND net1001 sg13g2_dlygate4sd3_1
Xhold222 _0034_ VPWR VGND net979 sg13g2_dlygate4sd3_1
Xhold233 _0236_ VPWR VGND net990 sg13g2_dlygate4sd3_1
X_4457_ net486 VPWR _1370_ VGND _1368_ _1369_ sg13g2_o21ai_1
Xhold266 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[4\] VPWR VGND net1023 sg13g2_dlygate4sd3_1
Xhold277 _1884_ VPWR VGND net1034 sg13g2_dlygate4sd3_1
Xhold255 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[9\] VPWR VGND
+ net1012 sg13g2_dlygate4sd3_1
X_6882__321 VPWR VGND net321 sg13g2_tiehi
Xhold299 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[5\] VPWR VGND net1056 sg13g2_dlygate4sd3_1
Xhold288 _0212_ VPWR VGND net1045 sg13g2_dlygate4sd3_1
X_4388_ VGND VPWR _1304_ _1309_ _0134_ _1310_ sg13g2_a21oi_1
X_6127_ _2753_ net1298 _2754_ VPWR VGND sg13g2_nor2b_1
X_6058_ _2686_ _2692_ _2693_ _2695_ VPWR VGND sg13g2_nor3_1
Xclkbuf_leaf_65_clk clknet_4_0_0_clk clknet_leaf_65_clk VPWR VGND sg13g2_buf_8
XFILLER_27_844 VPWR VGND sg13g2_fill_2
X_5009_ _1829_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[1\] _1828_
+ VPWR VGND sg13g2_nand2_1
XFILLER_6_748 VPWR VGND sg13g2_decap_8
XFILLER_2_921 VPWR VGND sg13g2_decap_8
X_6887__298 VPWR VGND net298 sg13g2_tiehi
XFILLER_2_998 VPWR VGND sg13g2_decap_8
X_6645__77 VPWR VGND net77 sg13g2_tiehi
XFILLER_37_619 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_56_clk clknet_4_10_0_clk clknet_leaf_56_clk VPWR VGND sg13g2_buf_8
XFILLER_18_822 VPWR VGND sg13g2_fill_1
XFILLER_17_343 VPWR VGND sg13g2_fill_1
XFILLER_29_192 VPWR VGND sg13g2_fill_2
X_6859__367 VPWR VGND net367 sg13g2_tiehi
XFILLER_33_858 VPWR VGND sg13g2_fill_1
XFILLER_32_379 VPWR VGND sg13g2_fill_2
XFILLER_9_520 VPWR VGND sg13g2_fill_2
X_3690_ _0743_ _0716_ _0742_ _0714_ _0713_ VPWR VGND sg13g2_a22oi_1
X_5360_ _2110_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[6\]
+ _2111_ VPWR VGND sg13g2_xor2_1
X_4311_ _1246_ _1249_ _1250_ VPWR VGND sg13g2_nor2_1
X_5291_ net1259 net528 _2053_ VPWR VGND sg13g2_xor2_1
X_4242_ _1190_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[1\]
+ _1189_ VPWR VGND sg13g2_xnor2_1
X_4173_ _1132_ net1574 _1130_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_47_clk clknet_4_8_0_clk clknet_leaf_47_clk VPWR VGND sg13g2_buf_8
X_6814_ net611 VGND VPWR _0423_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[9\]
+ clknet_leaf_59_clk sg13g2_dfrbpq_2
X_6745_ net680 VGND VPWR _0354_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[4\]\[3\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_1
XFILLER_11_519 VPWR VGND sg13g2_fill_2
X_3957_ net763 net1007 _0958_ VPWR VGND sg13g2_nor2_1
X_3888_ _0632_ _0904_ _0911_ VPWR VGND sg13g2_nor2_2
X_6676_ net46 VGND VPWR _0285_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[4\]
+ clknet_leaf_49_clk sg13g2_dfrbpq_2
X_5627_ VGND VPWR _2335_ _2336_ _2329_ _0598_ sg13g2_a21oi_2
X_5558_ VGND VPWR _2268_ _2274_ _2276_ net425 sg13g2_a21oi_1
X_4509_ VGND VPWR _1409_ _1413_ _0151_ _1414_ sg13g2_a21oi_1
X_5489_ _2212_ _2213_ _2218_ _2221_ VPWR VGND sg13g2_nor3_1
Xfanout521 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].z_sign net521
+ VPWR VGND sg13g2_buf_8
Xfanout510 net511 net510 VPWR VGND sg13g2_buf_8
Xfanout532 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].z_sign net532
+ VPWR VGND sg13g2_buf_2
Xfanout554 u_angle_cordic_12b_pmod.u_vga_top.pixel_clk_en net554 VPWR VGND sg13g2_buf_8
Xfanout543 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].z_sign net543
+ VPWR VGND sg13g2_buf_8
XFILLER_18_118 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_38_clk clknet_4_15_0_clk clknet_leaf_38_clk VPWR VGND sg13g2_buf_8
XFILLER_26_162 VPWR VGND sg13g2_fill_2
XFILLER_41_165 VPWR VGND sg13g2_fill_2
XFILLER_29_1004 VPWR VGND sg13g2_decap_8
XFILLER_2_795 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_29_clk clknet_4_9_0_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
X_4860_ _1705_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[1\]
+ _1704_ VPWR VGND sg13g2_xnor2_1
X_3811_ net552 net909 _0853_ VPWR VGND sg13g2_nor2_1
X_4791_ _1646_ _1647_ _1648_ VPWR VGND sg13g2_nor2b_1
X_6530_ net192 VGND VPWR _0139_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[6\]
+ clknet_leaf_32_clk sg13g2_dfrbpq_1
XFILLER_13_390 VPWR VGND sg13g2_fill_2
X_3742_ _0781_ _0783_ _0794_ _0795_ VPWR VGND sg13g2_nor3_1
X_6461_ net273 VGND VPWR _0070_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[0\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_2
X_3673_ _0644_ VPWR _0726_ VGND _0637_ _0638_ sg13g2_o21ai_1
X_5412_ net477 VPWR _2155_ VGND _2149_ _2154_ sg13g2_o21ai_1
X_6392_ net574 VGND VPWR _0001_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[0\].y_shr\[10\]
+ clknet_leaf_65_clk sg13g2_dfrbpq_2
X_5343_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[4\] VPWR _2096_
+ VGND _2087_ _2093_ sg13g2_o21ai_1
X_5274_ VGND VPWR net804 _2037_ _2039_ _2036_ sg13g2_a21oi_1
X_4225_ _1172_ _1175_ _1177_ VPWR VGND sg13g2_nor2_1
X_4156_ net534 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[6\] _1117_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_43_408 VPWR VGND sg13g2_fill_1
X_4087_ net420 _1065_ _1066_ _0076_ VPWR VGND sg13g2_nor3_1
XFILLER_11_338 VPWR VGND sg13g2_fill_1
X_4989_ VGND VPWR net1434 _1812_ _0232_ _1813_ sg13g2_a21oi_1
X_6728_ net697 VGND VPWR net812 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].z_sign
+ clknet_leaf_47_clk sg13g2_dfrbpq_1
X_6659_ net63 VGND VPWR net1164 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[6\]
+ clknet_leaf_50_clk sg13g2_dfrbpq_2
XFILLER_3_515 VPWR VGND sg13g2_fill_1
Xfanout373 _0991_ net373 VPWR VGND sg13g2_buf_8
Xfanout384 net385 net384 VPWR VGND sg13g2_buf_8
Xfanout395 _1843_ net395 VPWR VGND sg13g2_buf_8
XFILLER_4_1028 VPWR VGND sg13g2_fill_1
XFILLER_14_187 VPWR VGND sg13g2_fill_1
XFILLER_30_647 VPWR VGND sg13g2_fill_1
Xinput15 uio_in[5] net15 VPWR VGND sg13g2_buf_1
XFILLER_7_876 VPWR VGND sg13g2_decap_8
XFILLER_6_397 VPWR VGND sg13g2_fill_1
X_4010_ _1008_ _1007_ _1006_ VPWR VGND sg13g2_nand2b_1
XFILLER_19_961 VPWR VGND sg13g2_decap_8
XFILLER_46_780 VPWR VGND sg13g2_fill_2
X_5961_ _2619_ _2611_ _2613_ _2618_ VPWR VGND sg13g2_and3_1
X_4912_ net390 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[9\] _1749_
+ VPWR VGND sg13g2_xor2_1
X_5892_ _2559_ net1146 _2557_ VPWR VGND sg13g2_xnor2_1
XFILLER_33_452 VPWR VGND sg13g2_fill_1
X_4843_ _1690_ _1691_ _1689_ _1692_ VPWR VGND sg13g2_nand3_1
X_4774_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[9\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[8\]
+ _1634_ VPWR VGND sg13g2_nor2_1
X_6513_ net209 VGND VPWR _0122_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[1\]
+ clknet_leaf_38_clk sg13g2_dfrbpq_1
X_3725_ _0754_ net407 net409 _0778_ VPWR VGND sg13g2_a21o_1
Xclkbuf_leaf_9_clk clknet_4_3_0_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
X_6444_ net303 VGND VPWR _0053_ u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[10\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
X_3656_ VGND VPWR _0707_ _0708_ _0709_ _0702_ sg13g2_a21oi_1
X_6375_ VGND VPWR net1029 _2925_ _2926_ net375 sg13g2_a21oi_1
X_3587_ net546 u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[3\] u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[3\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[3\] net535 net544 _0640_
+ VPWR VGND sg13g2_mux4_1
X_5326_ _0556_ _2080_ _2081_ VPWR VGND sg13g2_nor2_1
X_5257_ _2028_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[6\]
+ net379 VPWR VGND sg13g2_xnor2_1
XFILLER_29_703 VPWR VGND sg13g2_fill_1
X_4208_ VGND VPWR _1155_ _1157_ _1163_ _1161_ sg13g2_a21oi_1
X_5188_ _1965_ VPWR _1968_ VGND _1961_ _1966_ sg13g2_o21ai_1
X_6410__360 VPWR VGND net360 sg13g2_tiehi
X_4139_ _1089_ _1091_ _1098_ _1101_ _1104_ VPWR VGND sg13g2_nor4_1
XFILLER_19_1003 VPWR VGND sg13g2_decap_8
XFILLER_25_975 VPWR VGND sg13g2_decap_8
XFILLER_11_113 VPWR VGND sg13g2_fill_2
XFILLER_12_636 VPWR VGND sg13g2_fill_1
XFILLER_40_945 VPWR VGND sg13g2_fill_1
Xheichips25_CORDIC_25 VPWR VGND uio_oe[1] sg13g2_tielo
XFILLER_4_846 VPWR VGND sg13g2_decap_8
Xheichips25_CORDIC_36 VPWR VGND uio_out[5] sg13g2_tielo
XFILLER_26_1007 VPWR VGND sg13g2_decap_8
XFILLER_47_83 VPWR VGND sg13g2_fill_2
XFILLER_47_61 VPWR VGND sg13g2_decap_8
XFILLER_47_599 VPWR VGND sg13g2_fill_1
XFILLER_16_942 VPWR VGND sg13g2_decap_8
XFILLER_28_780 VPWR VGND sg13g2_fill_2
XFILLER_15_441 VPWR VGND sg13g2_fill_1
XFILLER_30_466 VPWR VGND sg13g2_fill_1
X_3510_ VPWR _0580_ net1562 VGND sg13g2_inv_1
Xhold607 _1134_ VPWR VGND net1364 sg13g2_dlygate4sd3_1
X_4490_ VGND VPWR _1398_ _1397_ _1393_ sg13g2_or2_1
Xhold618 _1332_ VPWR VGND net1375 sg13g2_dlygate4sd3_1
Xhold629 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[11\] VPWR VGND net1386
+ sg13g2_dlygate4sd3_1
X_6160_ VPWR _2783_ _2782_ VGND sg13g2_inv_1
X_5111_ _1903_ net1485 _1901_ VPWR VGND sg13g2_xnor2_1
X_6091_ net424 net1372 _2723_ _0424_ VPWR VGND sg13g2_nor3_1
X_5042_ _1857_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[6\] _1843_
+ VPWR VGND sg13g2_nand2_1
XFILLER_38_577 VPWR VGND sg13g2_fill_1
XFILLER_19_780 VPWR VGND sg13g2_fill_1
X_5944_ _2604_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[10\] _2603_
+ VPWR VGND sg13g2_xnor2_1
X_5875_ _2542_ VPWR _2545_ VGND _2539_ _2543_ sg13g2_o21ai_1
XFILLER_22_923 VPWR VGND sg13g2_decap_8
X_4826_ _1671_ VPWR _1677_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[7\]
+ net391 sg13g2_o21ai_1
XFILLER_21_477 VPWR VGND sg13g2_fill_2
X_4757_ _1615_ _1618_ _1620_ VPWR VGND sg13g2_and2_1
XFILLER_49_1007 VPWR VGND sg13g2_decap_8
X_4688_ VGND VPWR net872 _1560_ _0183_ _1561_ sg13g2_a21oi_1
X_3708_ _0761_ _0749_ _0759_ VPWR VGND sg13g2_xnor2_1
X_7476_ net22 net19 VPWR VGND sg13g2_buf_1
X_6427_ net326 VGND VPWR _0036_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[5\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_2
X_3639_ _0690_ _0672_ _0692_ VPWR VGND sg13g2_xor2_1
XFILLER_1_805 VPWR VGND sg13g2_decap_8
X_6358_ net975 _2913_ _2915_ VPWR VGND sg13g2_and2_1
X_5309_ VPWR VGND _2066_ _2067_ _2056_ net415 _2068_ net1268 sg13g2_a221oi_1
X_6289_ net444 VPWR _2886_ VGND net555 _2881_ sg13g2_o21ai_1
XFILLER_44_536 VPWR VGND sg13g2_fill_2
XFILLER_13_923 VPWR VGND sg13g2_decap_8
XFILLER_0_871 VPWR VGND sg13g2_decap_8
Xhold4 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[0\] VPWR VGND net761
+ sg13g2_dlygate4sd3_1
XFILLER_16_750 VPWR VGND sg13g2_fill_1
X_3990_ _0991_ net448 _0986_ VPWR VGND sg13g2_nand2_1
X_5660_ _2362_ _2363_ _0353_ VPWR VGND sg13g2_nor2b_1
X_4611_ _1496_ net1165 _1494_ VPWR VGND sg13g2_xnor2_1
X_5591_ net474 VPWR _2305_ VGND _2300_ _2304_ sg13g2_o21ai_1
X_4542_ VGND VPWR _1439_ _1440_ _0157_ _1441_ sg13g2_a21oi_1
XFILLER_8_993 VPWR VGND sg13g2_decap_8
Xhold404 _0225_ VPWR VGND net1161 sg13g2_dlygate4sd3_1
Xhold415 _2263_ VPWR VGND net1172 sg13g2_dlygate4sd3_1
Xhold426 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[2\] VPWR
+ VGND net1183 sg13g2_dlygate4sd3_1
X_6869__347 VPWR VGND net347 sg13g2_tiehi
X_4473_ net487 VPWR _1383_ VGND _1377_ _1382_ sg13g2_o21ai_1
Xhold459 _0223_ VPWR VGND net1216 sg13g2_dlygate4sd3_1
Xhold437 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[11\] VPWR VGND net1194
+ sg13g2_dlygate4sd3_1
X_6212_ net426 _2824_ _2825_ _0443_ VPWR VGND sg13g2_nor3_1
Xhold448 _0368_ VPWR VGND net1205 sg13g2_dlygate4sd3_1
X_6143_ _2768_ net1406 _2766_ VPWR VGND sg13g2_xnor2_1
X_6074_ _2707_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[8\] _2709_
+ VPWR VGND sg13g2_xor2_1
X_5025_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].y_shr\[10\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].z_sign
+ _1834_ _1843_ VPWR VGND sg13g2_a21o_2
X_5927_ _2587_ _2582_ _2585_ _2589_ VPWR VGND sg13g2_a21o_1
XFILLER_10_915 VPWR VGND sg13g2_decap_8
X_5858_ _2531_ _2530_ _2525_ VPWR VGND sg13g2_nand2b_1
XFILLER_16_1028 VPWR VGND sg13g2_fill_1
X_5789_ net476 VPWR _2472_ VGND _2470_ _2471_ sg13g2_o21ai_1
X_4809_ _1659_ _1656_ _1662_ _1664_ VPWR VGND sg13g2_a21o_2
X_6852__384 VPWR VGND net568 sg13g2_tiehi
XFILLER_1_679 VPWR VGND sg13g2_decap_8
XFILLER_45_801 VPWR VGND sg13g2_fill_1
XFILLER_5_996 VPWR VGND sg13g2_decap_8
XFILLER_39_149 VPWR VGND sg13g2_fill_1
XFILLER_48_661 VPWR VGND sg13g2_fill_1
X_6830_ net595 VGND VPWR net1283 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[10\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_2
X_6761_ net664 VGND VPWR _0370_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[6\]
+ clknet_leaf_30_clk sg13g2_dfrbpq_1
XFILLER_35_377 VPWR VGND sg13g2_fill_2
XFILLER_16_580 VPWR VGND sg13g2_fill_1
X_5712_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[11\] net412 _2401_
+ _2409_ VPWR VGND sg13g2_a21o_1
X_6498__224 VPWR VGND net224 sg13g2_tiehi
X_3973_ _0963_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[10\] _0974_
+ VPWR VGND sg13g2_xor2_1
X_6692_ net747 VGND VPWR net1009 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[1\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_5643_ net1010 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[3\] _2349_
+ VPWR VGND sg13g2_nor2b_1
X_5574_ _2290_ net1384 _2287_ VPWR VGND sg13g2_xnor2_1
X_4525_ _1425_ _1427_ _1428_ VPWR VGND sg13g2_and2_1
Xhold201 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[13\] VPWR VGND net958
+ sg13g2_dlygate4sd3_1
Xhold223 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[2\] VPWR VGND
+ net980 sg13g2_dlygate4sd3_1
Xhold212 _0452_ VPWR VGND net969 sg13g2_dlygate4sd3_1
Xhold234 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[0\] VPWR
+ VGND net991 sg13g2_dlygate4sd3_1
Xhold267 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[1\] VPWR VGND net1024 sg13g2_dlygate4sd3_1
Xhold245 _0040_ VPWR VGND net1002 sg13g2_dlygate4sd3_1
Xhold278 _0262_ VPWR VGND net1035 sg13g2_dlygate4sd3_1
Xhold256 _0065_ VPWR VGND net1013 sg13g2_dlygate4sd3_1
X_4456_ VGND VPWR net1158 net386 _1369_ _1366_ sg13g2_a21oi_1
X_4387_ net502 VPWR _1310_ VGND _1304_ _1309_ sg13g2_o21ai_1
Xhold289 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[0\] VPWR VGND net1046
+ sg13g2_dlygate4sd3_1
X_6126_ _2752_ net1295 _2753_ VPWR VGND sg13g2_xor2_1
X_6057_ _2692_ VPWR _2694_ VGND _2686_ _2693_ sg13g2_o21ai_1
XFILLER_22_1021 VPWR VGND sg13g2_decap_8
X_5008_ _1828_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].y_shr\[1\]
+ _1827_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_322 VPWR VGND sg13g2_fill_1
XFILLER_27_856 VPWR VGND sg13g2_fill_1
XFILLER_26_399 VPWR VGND sg13g2_fill_1
XFILLER_6_727 VPWR VGND sg13g2_decap_8
XFILLER_2_900 VPWR VGND sg13g2_decap_8
Xhold790 _2761_ VPWR VGND net1547 sg13g2_dlygate4sd3_1
XFILLER_2_977 VPWR VGND sg13g2_decap_8
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk VPWR VGND sg13g2_buf_8
XFILLER_17_322 VPWR VGND sg13g2_fill_2
XFILLER_44_174 VPWR VGND sg13g2_fill_2
XFILLER_33_848 VPWR VGND sg13g2_fill_1
XFILLER_5_793 VPWR VGND sg13g2_decap_8
X_4310_ _1248_ VPWR _1249_ VGND _1241_ _1242_ sg13g2_o21ai_1
X_5290_ VGND VPWR _2048_ _2050_ _0294_ _2052_ sg13g2_a21oi_1
X_4241_ net531 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[0\]
+ _1189_ VPWR VGND sg13g2_nor2b_1
X_4172_ net534 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[9\] _1131_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_36_620 VPWR VGND sg13g2_fill_2
X_6813_ net612 VGND VPWR net1321 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[8\]
+ clknet_leaf_59_clk sg13g2_dfrbpq_1
X_6744_ net681 VGND VPWR _0353_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[4\]\[2\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3956_ _0942_ _0956_ _0957_ VPWR VGND sg13g2_nor2b_1
X_6675_ net47 VGND VPWR net1182 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[3\]
+ clknet_leaf_48_clk sg13g2_dfrbpq_2
X_3887_ _0535_ _0907_ _0910_ VPWR VGND sg13g2_and2_1
X_5626_ net412 _0598_ _2335_ VPWR VGND sg13g2_nor2_1
X_5557_ _2268_ _2274_ _2275_ VPWR VGND sg13g2_nor2_1
X_5488_ net430 _2219_ net1484 _0324_ VPWR VGND sg13g2_nor3_1
X_4508_ net498 VPWR _1414_ VGND _1409_ _1413_ sg13g2_o21ai_1
X_4439_ _1350_ VPWR _1355_ VGND _1343_ _1346_ sg13g2_o21ai_1
Xfanout511 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].z_sign net511
+ VPWR VGND sg13g2_buf_8
Xfanout522 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].z_sign net522
+ VPWR VGND sg13g2_buf_1
Xfanout533 net534 net533 VPWR VGND sg13g2_buf_8
Xfanout500 net505 net500 VPWR VGND sg13g2_buf_2
Xfanout555 net1043 net555 VPWR VGND sg13g2_buf_8
Xfanout544 net545 net544 VPWR VGND sg13g2_buf_8
X_6109_ _2738_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[2\] _2737_
+ VPWR VGND sg13g2_xnor2_1
X_6895__546 VPWR VGND net730 sg13g2_tiehi
X_6420__340 VPWR VGND net340 sg13g2_tiehi
XFILLER_2_774 VPWR VGND sg13g2_decap_8
X_6488__234 VPWR VGND net234 sg13g2_tiehi
XFILLER_1_295 VPWR VGND sg13g2_fill_2
XFILLER_46_984 VPWR VGND sg13g2_fill_1
XFILLER_33_601 VPWR VGND sg13g2_fill_2
X_6641__81 VPWR VGND net81 sg13g2_tiehi
XFILLER_33_634 VPWR VGND sg13g2_fill_1
X_4790_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[11\] _1645_ _0613_
+ _1647_ VPWR VGND sg13g2_nand3_1
X_3810_ VGND VPWR net552 _0851_ _0014_ net893 sg13g2_a21oi_1
XFILLER_14_892 VPWR VGND sg13g2_decap_8
X_3741_ _0793_ _0775_ _0794_ VPWR VGND sg13g2_xor2_1
X_6495__227 VPWR VGND net227 sg13g2_tiehi
X_6460_ net274 VGND VPWR _0069_ u_angle_cordic_12b_pmod.waveform_sel_reg\[1\] clknet_leaf_16_clk
+ sg13g2_dfrbpq_1
X_3672_ _0718_ _0638_ _0725_ VPWR VGND sg13g2_nor2b_1
X_6391_ net725 VGND VPWR _0000_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[0\].y_shr\[11\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_2
X_5411_ _2154_ net1304 _2152_ VPWR VGND sg13g2_xnor2_1
X_5342_ VPWR _2095_ _2094_ VGND sg13g2_inv_1
X_5273_ VGND VPWR net804 _2037_ _0291_ _2038_ sg13g2_a21oi_1
X_4224_ _1172_ _1175_ _1176_ VPWR VGND sg13g2_and2_1
X_4155_ net437 _1116_ _0095_ VPWR VGND sg13g2_nor2_1
X_4086_ _0531_ _1064_ _1066_ VPWR VGND sg13g2_nor2_2
XFILLER_23_166 VPWR VGND sg13g2_fill_1
X_6918__262 VPWR VGND net262 sg13g2_tiehi
X_4988_ net468 VPWR _1813_ VGND _1810_ _1812_ sg13g2_o21ai_1
X_3939_ _0940_ VPWR _0941_ VGND _0936_ _0937_ sg13g2_o21ai_1
X_6727_ net698 VGND VPWR net1126 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[10\]
+ clknet_leaf_47_clk sg13g2_dfrbpq_2
X_6658_ net64 VGND VPWR net1276 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[5\]
+ clknet_leaf_50_clk sg13g2_dfrbpq_1
X_5609_ _2318_ _2312_ _2316_ _2320_ VPWR VGND sg13g2_a21o_1
X_6589_ net133 VGND VPWR _0198_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[0\]
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
XFILLER_4_1007 VPWR VGND sg13g2_decap_8
Xfanout374 net375 net374 VPWR VGND sg13g2_buf_8
Xfanout396 _1842_ net396 VPWR VGND sg13g2_buf_8
Xfanout385 _1416_ net385 VPWR VGND sg13g2_buf_8
XFILLER_14_144 VPWR VGND sg13g2_fill_1
Xinput16 uio_in[6] net16 VPWR VGND sg13g2_buf_1
XFILLER_11_884 VPWR VGND sg13g2_decap_8
XFILLER_7_855 VPWR VGND sg13g2_decap_8
XFILLER_37_214 VPWR VGND sg13g2_fill_2
XFILLER_19_940 VPWR VGND sg13g2_decap_8
X_5960_ _2618_ net1530 _2616_ VPWR VGND sg13g2_xnor2_1
X_4911_ VGND VPWR _1744_ _1746_ _0219_ _1748_ sg13g2_a21oi_1
X_5891_ _2558_ net1146 _2557_ VPWR VGND sg13g2_nand2_1
XFILLER_34_987 VPWR VGND sg13g2_fill_1
X_4842_ net392 VPWR _1691_ VGND net1044 net1137 sg13g2_o21ai_1
X_4773_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[3\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[2\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[1\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[0\]
+ _1633_ VPWR VGND sg13g2_nor4_1
X_6512_ net210 VGND VPWR _0121_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[0\]
+ clknet_leaf_38_clk sg13g2_dfrbpq_1
X_3724_ _0777_ _0660_ _0754_ VPWR VGND sg13g2_nand2_1
X_6443_ net304 VGND VPWR _0052_ u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[9\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_1
X_3655_ _0701_ _0700_ _0708_ VPWR VGND sg13g2_xor2_1
X_6374_ net375 net917 _2925_ _0517_ VPWR VGND sg13g2_nor3_1
X_3586_ net547 u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[0\] u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[0\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[0\] net535 net545 _0639_
+ VPWR VGND sg13g2_mux4_1
X_5325_ _2080_ _0555_ _2079_ VPWR VGND sg13g2_xnor2_1
X_5256_ _0285_ net492 _2026_ _2027_ VPWR VGND sg13g2_and3_1
X_4207_ _1162_ _1155_ _1157_ _1161_ VPWR VGND sg13g2_and3_1
X_5187_ VGND VPWR _1961_ net1063 _0276_ _1967_ sg13g2_a21oi_1
X_6879__327 VPWR VGND net327 sg13g2_tiehi
XFILLER_28_236 VPWR VGND sg13g2_fill_2
X_4138_ net437 _1102_ net1151 _0091_ VPWR VGND sg13g2_nor3_1
X_4069_ _1054_ _1053_ net840 VPWR VGND sg13g2_nand2b_1
XFILLER_25_954 VPWR VGND sg13g2_decap_8
X_6478__244 VPWR VGND net244 sg13g2_tiehi
XFILLER_4_825 VPWR VGND sg13g2_decap_8
Xheichips25_CORDIC_26 VPWR VGND uio_oe[2] sg13g2_tielo
Xheichips25_CORDIC_37 VPWR VGND uio_out[6] sg13g2_tielo
XFILLER_19_203 VPWR VGND sg13g2_fill_1
X_6485__237 VPWR VGND net237 sg13g2_tiehi
XFILLER_16_921 VPWR VGND sg13g2_decap_8
XFILLER_34_217 VPWR VGND sg13g2_fill_2
XFILLER_43_740 VPWR VGND sg13g2_fill_2
XFILLER_16_998 VPWR VGND sg13g2_decap_8
Xhold608 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[1\] VPWR VGND net1365
+ sg13g2_dlygate4sd3_1
Xhold619 _0137_ VPWR VGND net1376 sg13g2_dlygate4sd3_1
X_6090_ VGND VPWR _2714_ _2717_ _2723_ _2721_ sg13g2_a21oi_1
X_5110_ _1902_ net1485 _1901_ VPWR VGND sg13g2_nand2_1
X_5041_ _1855_ VPWR _1856_ VGND _1850_ _1853_ sg13g2_o21ai_1
X_5943_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[9\] net413 _2597_
+ _2603_ VPWR VGND sg13g2_a21o_1
X_5874_ VGND VPWR _2539_ net1423 _0386_ _2544_ sg13g2_a21oi_1
XFILLER_22_979 VPWR VGND sg13g2_decap_8
X_4825_ VGND VPWR _1674_ _1675_ _0205_ _1676_ sg13g2_a21oi_1
X_4756_ _1615_ _1618_ _1619_ VPWR VGND sg13g2_nor2_1
X_4687_ net488 VPWR _1561_ VGND net872 _1560_ sg13g2_o21ai_1
X_7475_ net21 net18 VPWR VGND sg13g2_buf_1
X_3707_ _0760_ _0759_ _0749_ VPWR VGND sg13g2_nand2b_1
X_6426_ net328 VGND VPWR _0035_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[4\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_2
X_3638_ _0672_ _0690_ _0691_ VPWR VGND sg13g2_nor2_1
X_3569_ u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[6\] u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[5\]
+ u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[4\] _0628_ VPWR VGND sg13g2_nor3_1
X_6357_ net374 _2913_ net881 _0511_ VPWR VGND sg13g2_nor3_1
X_5308_ _2067_ _2059_ _2057_ VPWR VGND sg13g2_nand2b_1
X_6288_ _0465_ net444 _2884_ _2885_ VPWR VGND sg13g2_and3_1
X_5239_ net430 net1539 _2013_ _0282_ VPWR VGND sg13g2_nor3_1
XFILLER_29_589 VPWR VGND sg13g2_fill_1
XFILLER_13_902 VPWR VGND sg13g2_decap_8
XFILLER_25_773 VPWR VGND sg13g2_fill_1
XFILLER_40_710 VPWR VGND sg13g2_fill_2
XFILLER_12_434 VPWR VGND sg13g2_fill_1
XFILLER_33_20 VPWR VGND sg13g2_fill_1
XFILLER_9_939 VPWR VGND sg13g2_decap_8
XFILLER_12_467 VPWR VGND sg13g2_fill_2
XFILLER_13_979 VPWR VGND sg13g2_decap_8
XFILLER_8_449 VPWR VGND sg13g2_fill_1
XFILLER_4_699 VPWR VGND sg13g2_decap_8
XFILLER_0_850 VPWR VGND sg13g2_decap_8
Xhold5 _0440_ VPWR VGND net762 sg13g2_dlygate4sd3_1
X_4610_ _1495_ net1165 _1494_ VPWR VGND sg13g2_nand2_1
X_5590_ _2304_ _0596_ _2302_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_798 VPWR VGND sg13g2_fill_2
X_4541_ net498 VPWR _1441_ VGND _1439_ _1440_ sg13g2_o21ai_1
XFILLER_8_972 VPWR VGND sg13g2_decap_8
Xhold416 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[8\] VPWR VGND net1173
+ sg13g2_dlygate4sd3_1
Xhold405 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[6\] VPWR VGND net1162
+ sg13g2_dlygate4sd3_1
Xhold427 _0104_ VPWR VGND net1184 sg13g2_dlygate4sd3_1
X_4472_ _1382_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[1\] _1380_
+ VPWR VGND sg13g2_xnor2_1
Xhold438 _0349_ VPWR VGND net1195 sg13g2_dlygate4sd3_1
X_6211_ VGND VPWR _2819_ _2821_ _2825_ _2823_ sg13g2_a21oi_1
Xhold449 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[3\] VPWR VGND net1206
+ sg13g2_dlygate4sd3_1
X_6142_ _2767_ net1406 _2766_ VPWR VGND sg13g2_nand2_1
X_6073_ _2708_ net1497 _2707_ VPWR VGND sg13g2_nand2b_1
X_5024_ VGND VPWR _1834_ _1842_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].y_shr\[10\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].z_sign sg13g2_a21oi_2
X_5926_ VGND VPWR _2582_ _2587_ _0394_ _2588_ sg13g2_a21oi_1
XFILLER_34_581 VPWR VGND sg13g2_fill_2
X_5857_ _2530_ _2529_ _2528_ VPWR VGND sg13g2_nand2b_1
XFILLER_6_909 VPWR VGND sg13g2_decap_8
X_5788_ net826 net520 _2471_ VPWR VGND sg13g2_xor2_1
X_4808_ _1659_ _1662_ _1656_ _1663_ VPWR VGND sg13g2_nand3_1
X_4739_ _1605_ _1603_ _1604_ VPWR VGND sg13g2_nand2_1
X_6475__247 VPWR VGND net247 sg13g2_tiehi
X_6409_ net362 VGND VPWR net871 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[7\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
X_6451__291 VPWR VGND net291 sg13g2_tiehi
XFILLER_1_636 VPWR VGND sg13g2_fill_1
XFILLER_1_658 VPWR VGND sg13g2_decap_8
X_6657__65 VPWR VGND net65 sg13g2_tiehi
XFILLER_29_342 VPWR VGND sg13g2_fill_1
XFILLER_45_824 VPWR VGND sg13g2_fill_1
XFILLER_32_518 VPWR VGND sg13g2_decap_4
XFILLER_13_721 VPWR VGND sg13g2_fill_1
XFILLER_12_297 VPWR VGND sg13g2_fill_1
XFILLER_5_975 VPWR VGND sg13g2_decap_8
XFILLER_5_57 VPWR VGND sg13g2_fill_1
X_6430__320 VPWR VGND net320 sg13g2_tiehi
XFILLER_39_106 VPWR VGND sg13g2_fill_2
X_6799__442 VPWR VGND net626 sg13g2_tiehi
X_6760_ net665 VGND VPWR net1085 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[5\]
+ clknet_leaf_29_clk sg13g2_dfrbpq_1
X_5711_ VGND VPWR _2400_ _2405_ _2408_ _2403_ sg13g2_a21oi_1
X_3972_ _0973_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[9\] _0955_
+ VPWR VGND sg13g2_xnor2_1
X_6691_ net748 VGND VPWR net972 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[0\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_5642_ VGND VPWR _2346_ _2347_ _0350_ _2348_ sg13g2_a21oi_1
X_6398__381 VPWR VGND net565 sg13g2_tiehi
X_5573_ VPWR _2289_ _2288_ VGND sg13g2_inv_1
X_4524_ _1422_ _1426_ _1427_ VPWR VGND sg13g2_nor2_1
Xhold202 _2920_ VPWR VGND net959 sg13g2_dlygate4sd3_1
Xhold213 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[0\] VPWR VGND net970
+ sg13g2_dlygate4sd3_1
Xhold235 _0109_ VPWR VGND net992 sg13g2_dlygate4sd3_1
Xhold224 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[12\] VPWR VGND net981
+ sg13g2_dlygate4sd3_1
XFILLER_49_19 VPWR VGND sg13g2_decap_8
Xhold268 _0032_ VPWR VGND net1025 sg13g2_dlygate4sd3_1
Xhold257 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[0\] VPWR VGND net1014
+ sg13g2_dlygate4sd3_1
Xhold246 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[4\] VPWR VGND net1003 sg13g2_dlygate4sd3_1
X_4455_ _1368_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[4\]
+ net386 VPWR VGND sg13g2_xnor2_1
Xhold279 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[10\] VPWR VGND net1036
+ sg13g2_dlygate4sd3_1
X_4386_ _1309_ net1097 _1307_ VPWR VGND sg13g2_xnor2_1
X_6125_ VGND VPWR _0619_ _2743_ _2752_ net507 sg13g2_a21oi_1
XFILLER_22_1000 VPWR VGND sg13g2_decap_8
X_6056_ VPWR VGND net1209 _2679_ _2685_ _2676_ _2693_ _2681_ sg13g2_a221oi_1
X_6654__68 VPWR VGND net68 sg13g2_tiehi
XFILLER_27_846 VPWR VGND sg13g2_fill_1
X_5007_ _1827_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].y_shr\[0\]
+ _0617_ VPWR VGND sg13g2_nand2_1
X_6407__366 VPWR VGND net366 sg13g2_tiehi
XFILLER_42_849 VPWR VGND sg13g2_fill_2
X_5909_ VGND VPWR _2568_ net1510 _0392_ _2573_ sg13g2_a21oi_1
X_6889_ net294 VGND VPWR _0498_ u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[9\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_1
Xhold791 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[10\] VPWR VGND net1548
+ sg13g2_dlygate4sd3_1
Xhold780 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[7\] VPWR VGND net1537
+ sg13g2_dlygate4sd3_1
XFILLER_2_956 VPWR VGND sg13g2_decap_8
XFILLER_7_1016 VPWR VGND sg13g2_decap_8
XFILLER_7_1027 VPWR VGND sg13g2_fill_2
XFILLER_36_109 VPWR VGND sg13g2_fill_1
XFILLER_29_194 VPWR VGND sg13g2_fill_1
XFILLER_9_511 VPWR VGND sg13g2_fill_1
XFILLER_9_566 VPWR VGND sg13g2_fill_2
XFILLER_5_772 VPWR VGND sg13g2_decap_8
XFILLER_4_282 VPWR VGND sg13g2_fill_2
X_4240_ net963 _1187_ _0108_ VPWR VGND sg13g2_nor2b_1
X_4171_ _1123_ VPWR _1130_ VGND net534 _0586_ sg13g2_o21ai_1
X_6812_ net613 VGND VPWR _0421_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[7\]
+ clknet_leaf_59_clk sg13g2_dfrbpq_2
X_6743_ net682 VGND VPWR net1241 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[4\]\[1\]
+ clknet_leaf_53_clk sg13g2_dfrbpq_1
X_3955_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[2\] VPWR _0956_
+ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt_sum\[5\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[1\]
+ sg13g2_o21ai_1
X_6674_ net48 VGND VPWR _0283_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[2\]
+ clknet_leaf_46_clk sg13g2_dfrbpq_2
X_3886_ _0906_ VPWR _0033_ VGND _0908_ _0909_ sg13g2_o21ai_1
X_5625_ _2332_ _2328_ _2331_ _2334_ VPWR VGND sg13g2_a21o_1
X_5556_ _2272_ _2273_ _2274_ VPWR VGND sg13g2_nor2b_1
X_5487_ VGND VPWR _2211_ _2217_ _2220_ _2218_ sg13g2_a21oi_1
X_4507_ _1411_ net1461 _1413_ VPWR VGND sg13g2_xor2_1
X_4438_ _1354_ net1472 net386 VPWR VGND sg13g2_xnor2_1
Xfanout512 net514 net512 VPWR VGND sg13g2_buf_8
Xfanout523 net525 net523 VPWR VGND sg13g2_buf_8
Xfanout501 net504 net501 VPWR VGND sg13g2_buf_8
Xfanout534 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].z_sign net534
+ VPWR VGND sg13g2_buf_8
X_4369_ _1294_ VPWR _1296_ VGND net541 _0607_ sg13g2_o21ai_1
Xfanout545 u_angle_cordic_12b_pmod.waveform_sel_reg\[1\] net545 VPWR VGND sg13g2_buf_2
X_6108_ net507 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[1\] _2737_
+ VPWR VGND sg13g2_nor2b_1
X_6039_ _2677_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[4\]
+ _2678_ VPWR VGND sg13g2_xor2_1
XFILLER_41_64 VPWR VGND sg13g2_fill_2
X_6789__452 VPWR VGND net636 sg13g2_tiehi
XFILLER_9_0 VPWR VGND sg13g2_fill_2
XFILLER_2_753 VPWR VGND sg13g2_decap_8
X_6796__445 VPWR VGND net629 sg13g2_tiehi
XFILLER_32_156 VPWR VGND sg13g2_fill_1
X_3740_ _0791_ _0789_ _0793_ VPWR VGND sg13g2_xor2_1
X_3671_ _0638_ _0640_ _0724_ VPWR VGND sg13g2_and2_1
X_6390_ VGND VPWR _2870_ _2887_ _0476_ _2894_ sg13g2_a21oi_1
X_5410_ _2153_ net1304 _2152_ VPWR VGND sg13g2_nand2_1
X_5341_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[4\] _2087_
+ _2093_ _2094_ VPWR VGND sg13g2_nor3_2
X_5272_ net487 VPWR _2038_ VGND net804 _2037_ sg13g2_o21ai_1
X_4223_ _1173_ _1174_ _1175_ VPWR VGND sg13g2_and2_1
X_4154_ _1116_ net1103 net1106 VPWR VGND sg13g2_xnor2_1
X_4085_ _0531_ _1064_ _1065_ VPWR VGND sg13g2_and2_1
X_6726_ net699 VGND VPWR _0335_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[9\]
+ clknet_leaf_47_clk sg13g2_dfrbpq_2
X_4987_ _1812_ net1421 net398 VPWR VGND sg13g2_xnor2_1
X_3938_ VGND VPWR _0940_ _0938_ net551 sg13g2_or2_1
X_3869_ net441 VPWR _0896_ VGND _0538_ _0894_ sg13g2_o21ai_1
X_6657_ net65 VGND VPWR _0266_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[4\]
+ clknet_leaf_49_clk sg13g2_dfrbpq_1
X_6588_ net134 VGND VPWR net1143 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].z_sign
+ clknet_leaf_24_clk sg13g2_dfrbpq_2
X_5608_ VGND VPWR _2312_ _2318_ _0345_ _2319_ sg13g2_a21oi_1
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk VPWR VGND sg13g2_buf_8
X_5539_ net1124 _0553_ _2260_ _2261_ VPWR VGND sg13g2_a21o_1
Xfanout375 _0989_ net375 VPWR VGND sg13g2_buf_8
Xfanout397 net398 net397 VPWR VGND sg13g2_buf_8
Xfanout386 net387 net386 VPWR VGND sg13g2_buf_8
XFILLER_46_248 VPWR VGND sg13g2_fill_1
X_6903__554 VPWR VGND net738 sg13g2_tiehi
XFILLER_28_985 VPWR VGND sg13g2_decap_8
XFILLER_36_86 VPWR VGND sg13g2_fill_1
XFILLER_11_841 VPWR VGND sg13g2_fill_2
XFILLER_7_834 VPWR VGND sg13g2_decap_8
XFILLER_6_377 VPWR VGND sg13g2_fill_1
XFILLER_46_760 VPWR VGND sg13g2_fill_2
XFILLER_18_440 VPWR VGND sg13g2_fill_2
X_4910_ _1748_ net484 _1747_ VPWR VGND sg13g2_nand2_1
X_5890_ _2557_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[3\] _2556_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_19_996 VPWR VGND sg13g2_decap_8
X_4841_ _1690_ _1683_ _1685_ VPWR VGND sg13g2_nand2_1
X_4772_ net536 VPWR _1632_ VGND _1629_ _1631_ sg13g2_o21ai_1
XFILLER_14_690 VPWR VGND sg13g2_fill_2
X_3723_ _0753_ net404 _0776_ VPWR VGND sg13g2_xor2_1
X_6511_ net211 VGND VPWR net1200 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[12\]
+ clknet_leaf_44_clk sg13g2_dfrbpq_2
X_6442_ net305 VGND VPWR _0051_ u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[8\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_1
X_3654_ VPWR _0707_ _0706_ VGND sg13g2_inv_1
X_3585_ net546 u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[2\] u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[2\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[2\] net535 net544 _0638_
+ VPWR VGND sg13g2_mux4_1
X_6373_ _2925_ net854 net916 _2921_ VPWR VGND sg13g2_and3_1
X_5324_ net418 VPWR _2079_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[0\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[1\] sg13g2_o21ai_1
X_5255_ _2025_ _2024_ _2023_ _2027_ VPWR VGND sg13g2_a21o_1
X_4206_ _1161_ net1208 net382 VPWR VGND sg13g2_xnor2_1
X_5186_ net494 VPWR _1967_ VGND _1961_ _1966_ sg13g2_o21ai_1
X_4137_ VGND VPWR _1097_ _1099_ _1103_ net1150 sg13g2_a21oi_1
X_4068_ _0992_ net378 net879 _0070_ VPWR VGND sg13g2_mux2_1
X_6779__462 VPWR VGND net646 sg13g2_tiehi
XFILLER_7_108 VPWR VGND sg13g2_fill_1
X_6709_ net716 VGND VPWR _0318_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[0\]
+ clknet_leaf_55_clk sg13g2_dfrbpq_2
XFILLER_4_804 VPWR VGND sg13g2_decap_8
XFILLER_3_336 VPWR VGND sg13g2_fill_1
Xheichips25_CORDIC_38 VPWR VGND uo_out[2] sg13g2_tielo
Xheichips25_CORDIC_27 VPWR VGND uio_oe[3] sg13g2_tielo
X_6786__455 VPWR VGND net639 sg13g2_tiehi
XFILLER_47_30 VPWR VGND sg13g2_fill_1
XFILLER_47_85 VPWR VGND sg13g2_fill_1
XFILLER_16_900 VPWR VGND sg13g2_decap_8
XFILLER_16_977 VPWR VGND sg13g2_decap_8
XFILLER_31_936 VPWR VGND sg13g2_fill_2
X_6793__448 VPWR VGND net632 sg13g2_tiehi
XFILLER_11_682 VPWR VGND sg13g2_fill_2
Xhold609 _0199_ VPWR VGND net1366 sg13g2_dlygate4sd3_1
XFILLER_3_892 VPWR VGND sg13g2_decap_8
X_5040_ net395 VPWR _1855_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[4\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[5\] sg13g2_o21ai_1
X_6908__284 VPWR VGND net284 sg13g2_tiehi
X_5942_ VGND VPWR _2596_ _2600_ _2602_ _2599_ sg13g2_a21oi_1
X_5873_ net459 VPWR _2544_ VGND _2539_ _2543_ sg13g2_o21ai_1
XFILLER_22_958 VPWR VGND sg13g2_decap_8
X_4824_ net468 VPWR _1676_ VGND _1674_ _1675_ sg13g2_o21ai_1
X_4755_ _1618_ _1616_ _1617_ VPWR VGND sg13g2_nand2_1
X_3706_ _0759_ _0751_ _0758_ VPWR VGND sg13g2_xnor2_1
X_7474_ pwm_data net17 VPWR VGND sg13g2_buf_1
X_4686_ _1559_ _1554_ _1557_ _1560_ VPWR VGND sg13g2_mux2_1
X_6425_ net330 VGND VPWR net979 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[3\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_2
X_3637_ _0690_ net406 _0688_ VPWR VGND sg13g2_xnor2_1
X_3568_ _0627_ _0538_ u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[9\] VPWR VGND sg13g2_nand2_1
X_6356_ VGND VPWR net847 _2910_ _2914_ net880 sg13g2_a21oi_1
X_5307_ _2060_ _2063_ _2066_ VPWR VGND sg13g2_nor2_1
X_6287_ _2885_ net402 _2883_ VPWR VGND sg13g2_nand2b_1
X_3499_ VPWR _0569_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[8\] VGND
+ sg13g2_inv_1
X_5238_ _2011_ _2005_ _2013_ VPWR VGND sg13g2_nor2b_1
X_5169_ _1951_ VPWR _1953_ VGND _0571_ net380 sg13g2_o21ai_1
XFILLER_44_538 VPWR VGND sg13g2_fill_1
XFILLER_44_549 VPWR VGND sg13g2_fill_2
XFILLER_25_741 VPWR VGND sg13g2_fill_2
XFILLER_24_251 VPWR VGND sg13g2_fill_1
XFILLER_9_918 VPWR VGND sg13g2_decap_8
XFILLER_13_958 VPWR VGND sg13g2_decap_8
X_6491__231 VPWR VGND net231 sg13g2_tiehi
X_6417__346 VPWR VGND net346 sg13g2_tiehi
XFILLER_4_645 VPWR VGND sg13g2_fill_1
Xhold6 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[0\] VPWR VGND net763
+ sg13g2_dlygate4sd3_1
XFILLER_12_991 VPWR VGND sg13g2_decap_8
X_4540_ VGND VPWR net1169 net384 _1440_ _1437_ sg13g2_a21oi_1
XFILLER_8_951 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_10_clk clknet_4_9_0_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
Xhold417 _0220_ VPWR VGND net1174 sg13g2_dlygate4sd3_1
Xhold406 _1926_ VPWR VGND net1163 sg13g2_dlygate4sd3_1
X_4471_ _1381_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[1\] _1380_
+ VPWR VGND sg13g2_nand2_1
Xhold439 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].y_shr\[1\] VPWR
+ VGND net1196 sg13g2_dlygate4sd3_1
X_6210_ _2824_ _2819_ _2821_ _2823_ VPWR VGND sg13g2_and3_1
Xhold428 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[9\] VPWR VGND net1185
+ sg13g2_dlygate4sd3_1
X_6141_ _2766_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[6\] _2765_
+ VPWR VGND sg13g2_xnor2_1
X_6769__472 VPWR VGND net656 sg13g2_tiehi
X_6072_ _2707_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[8\]
+ _2706_ VPWR VGND sg13g2_xnor2_1
X_5023_ VGND VPWR _1832_ _1838_ _1841_ _1837_ sg13g2_a21oi_1
XFILLER_0_1011 VPWR VGND sg13g2_decap_8
X_5925_ net458 VPWR _2588_ VGND _2582_ _2587_ sg13g2_o21ai_1
X_5856_ _2529_ _0580_ _2527_ VPWR VGND sg13g2_nand2_1
X_6776__465 VPWR VGND net649 sg13g2_tiehi
XFILLER_16_1019 VPWR VGND sg13g2_decap_8
X_4807_ _1662_ net1237 net392 VPWR VGND sg13g2_xnor2_1
X_5787_ VGND VPWR _0592_ net1127 _2470_ _2469_ sg13g2_a21oi_1
X_4738_ VGND VPWR _1604_ net400 net1458 sg13g2_or2_1
X_4669_ net485 VPWR _1546_ VGND _1544_ _1545_ sg13g2_o21ai_1
X_6408_ net364 VGND VPWR net868 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[6\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_1
XFILLER_1_626 VPWR VGND sg13g2_fill_1
X_6339_ net926 _2901_ _2903_ VPWR VGND sg13g2_and2_1
X_6783__458 VPWR VGND net642 sg13g2_tiehi
XFILLER_44_346 VPWR VGND sg13g2_fill_1
XFILLER_32_508 VPWR VGND sg13g2_fill_2
XFILLER_40_530 VPWR VGND sg13g2_fill_1
XFILLER_8_203 VPWR VGND sg13g2_fill_2
XFILLER_5_954 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_59_clk clknet_4_3_0_clk clknet_leaf_59_clk VPWR VGND sg13g2_buf_8
XFILLER_36_803 VPWR VGND sg13g2_fill_2
XFILLER_35_313 VPWR VGND sg13g2_fill_2
X_3971_ _0966_ _0970_ _0961_ _0972_ VPWR VGND _0971_ sg13g2_nand4_1
X_5710_ net431 net1520 _2407_ _0359_ VPWR VGND sg13g2_nor3_1
X_6690_ net749 VGND VPWR net838 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].z_sign
+ clknet_leaf_44_clk sg13g2_dfrbpq_2
X_5641_ net476 VPWR _2348_ VGND _2346_ _2347_ sg13g2_o21ai_1
X_5572_ _2288_ net1384 _2287_ VPWR VGND sg13g2_nand2_1
X_4523_ VPWR VGND _1415_ _1417_ _1418_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[7\]
+ _1426_ net384 sg13g2_a221oi_1
Xhold214 _2072_ VPWR VGND net971 sg13g2_dlygate4sd3_1
Xhold203 _0514_ VPWR VGND net960 sg13g2_dlygate4sd3_1
Xhold225 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[10\] VPWR VGND
+ net982 sg13g2_dlygate4sd3_1
Xhold269 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[2\] VPWR VGND net1026
+ sg13g2_dlygate4sd3_1
X_4454_ VGND VPWR _1363_ _1365_ _0143_ _1367_ sg13g2_a21oi_1
Xhold258 _2474_ VPWR VGND net1015 sg13g2_dlygate4sd3_1
Xhold247 _0913_ VPWR VGND net1004 sg13g2_dlygate4sd3_1
Xhold236 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[0\] VPWR VGND net993
+ sg13g2_dlygate4sd3_1
X_4385_ _1308_ net1097 _1307_ VPWR VGND sg13g2_nand2_1
X_6124_ _2747_ _2742_ _2746_ _2751_ VPWR VGND sg13g2_a21o_1
X_6055_ _2692_ net1522 _2690_ VPWR VGND sg13g2_xnor2_1
X_5006_ net989 _1825_ _0236_ VPWR VGND sg13g2_nor2b_1
XFILLER_26_313 VPWR VGND sg13g2_fill_1
XFILLER_27_825 VPWR VGND sg13g2_fill_1
X_6481__241 VPWR VGND net241 sg13g2_tiehi
X_5908_ net457 VPWR _2573_ VGND _2568_ _2572_ sg13g2_o21ai_1
X_6888_ net296 VGND VPWR _0497_ u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[8\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_1
X_5839_ _2513_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[6\]
+ _2514_ VPWR VGND sg13g2_xor2_1
XFILLER_2_935 VPWR VGND sg13g2_decap_8
Xhold781 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[1\] VPWR
+ VGND net1538 sg13g2_dlygate4sd3_1
Xhold770 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[10\] VPWR VGND net1527
+ sg13g2_dlygate4sd3_1
Xhold792 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[7\] VPWR
+ VGND net1549 sg13g2_dlygate4sd3_1
XFILLER_17_313 VPWR VGND sg13g2_fill_2
XFILLER_17_324 VPWR VGND sg13g2_fill_1
X_6597__125 VPWR VGND net125 sg13g2_tiehi
X_6759__482 VPWR VGND net666 sg13g2_tiehi
XFILLER_9_556 VPWR VGND sg13g2_fill_1
XFILLER_5_751 VPWR VGND sg13g2_decap_8
XFILLER_45_1023 VPWR VGND sg13g2_fill_2
X_4170_ _1126_ _1122_ _1125_ _1129_ VPWR VGND sg13g2_a21o_1
X_6766__475 VPWR VGND net659 sg13g2_tiehi
XFILLER_36_622 VPWR VGND sg13g2_fill_1
X_6811_ net614 VGND VPWR _0420_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[6\]
+ clknet_leaf_59_clk sg13g2_dfrbpq_2
X_6697__558 VPWR VGND net742 sg13g2_tiehi
XFILLER_36_699 VPWR VGND sg13g2_fill_1
X_6742_ net683 VGND VPWR _0351_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[4\]\[0\]
+ clknet_leaf_54_clk sg13g2_dfrbpq_1
X_3954_ _0955_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[4\] _0943_
+ VPWR VGND sg13g2_xnor2_1
X_6673_ net49 VGND VPWR net1540 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[1\]
+ clknet_leaf_46_clk sg13g2_dfrbpq_2
X_3885_ _0909_ net443 _0901_ VPWR VGND sg13g2_nand2_1
X_6773__468 VPWR VGND net652 sg13g2_tiehi
X_5624_ VGND VPWR _2328_ _2332_ _0347_ _2333_ sg13g2_a21oi_1
X_5555_ _2273_ _0593_ _2271_ VPWR VGND sg13g2_nand2_1
X_5486_ _2219_ _2211_ _2217_ _2218_ VPWR VGND sg13g2_and3_1
X_4506_ _1412_ net1461 _1411_ VPWR VGND sg13g2_nand2b_1
X_4437_ _1353_ net1472 net386 VPWR VGND sg13g2_nand2_1
Xfanout513 net514 net513 VPWR VGND sg13g2_buf_8
Xfanout524 net525 net524 VPWR VGND sg13g2_buf_2
Xfanout502 net504 net502 VPWR VGND sg13g2_buf_8
Xfanout546 net547 net546 VPWR VGND sg13g2_buf_8
X_6107_ net424 net966 _0427_ VPWR VGND sg13g2_nor2_1
Xfanout535 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp\[0\] net535
+ VPWR VGND sg13g2_buf_2
X_4368_ VGND VPWR _1292_ _1293_ _0129_ _1295_ sg13g2_a21oi_1
X_4299_ _1235_ _1238_ _1239_ _1240_ VPWR VGND sg13g2_or3_1
X_6038_ VGND VPWR _0620_ _2668_ _2677_ net507 sg13g2_a21oi_1
XFILLER_26_187 VPWR VGND sg13g2_fill_2
X_6650__72 VPWR VGND net72 sg13g2_tiehi
XFILLER_2_732 VPWR VGND sg13g2_decap_8
XFILLER_29_1018 VPWR VGND sg13g2_decap_8
XFILLER_1_220 VPWR VGND sg13g2_fill_2
XFILLER_17_132 VPWR VGND sg13g2_fill_1
XFILLER_14_850 VPWR VGND sg13g2_fill_1
X_3670_ _0717_ _0722_ _0723_ VPWR VGND sg13g2_nor2_1
X_5340_ net521 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[3\]
+ _2093_ VPWR VGND sg13g2_nor2b_1
X_5271_ _2037_ net528 net862 VPWR VGND sg13g2_xnor2_1
X_4222_ net383 VPWR _1174_ VGND net1183 net1559 sg13g2_o21ai_1
X_4153_ net1103 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[6\] _1115_
+ VPWR VGND sg13g2_nor2b_1
X_4084_ _0075_ net445 _1063_ _1064_ VPWR VGND sg13g2_and3_1
XFILLER_36_463 VPWR VGND sg13g2_fill_2
X_4986_ _1811_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[8\] net397
+ VPWR VGND sg13g2_nand2_1
X_6725_ net700 VGND VPWR _0334_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[8\]
+ clknet_leaf_47_clk sg13g2_dfrbpq_2
X_3937_ _0939_ net918 net548 VPWR VGND sg13g2_nand2b_1
X_3868_ net888 _0895_ _0029_ VPWR VGND sg13g2_nor2_1
X_6656_ net66 VGND VPWR _0265_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[3\]
+ clknet_leaf_48_clk sg13g2_dfrbpq_1
X_6587_ net135 VGND VPWR net1400 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[12\]
+ clknet_leaf_34_clk sg13g2_dfrbpq_2
X_3799_ _0845_ _0826_ net1066 _0010_ VPWR VGND sg13g2_a21o_1
X_5607_ net475 VPWR _2319_ VGND _2312_ _2318_ sg13g2_o21ai_1
X_5538_ net432 _2259_ _2260_ _0334_ VPWR VGND sg13g2_nor3_1
X_5469_ _2205_ _2199_ _2203_ VPWR VGND sg13g2_nand2b_1
X_6587__135 VPWR VGND net135 sg13g2_tiehi
X_6749__492 VPWR VGND net676 sg13g2_tiehi
Xfanout376 net377 net376 VPWR VGND sg13g2_buf_8
Xfanout398 net399 net398 VPWR VGND sg13g2_buf_8
Xfanout387 _1342_ net387 VPWR VGND sg13g2_buf_8
X_6448__297 VPWR VGND net297 sg13g2_tiehi
XFILLER_36_65 VPWR VGND sg13g2_fill_1
X_6594__128 VPWR VGND net128 sg13g2_tiehi
X_6756__485 VPWR VGND net669 sg13g2_tiehi
XFILLER_7_813 VPWR VGND sg13g2_decap_8
X_6687__568 VPWR VGND net752 sg13g2_tiehi
XFILLER_35_8 VPWR VGND sg13g2_fill_1
X_6763__478 VPWR VGND net662 sg13g2_tiehi
X_6427__326 VPWR VGND net326 sg13g2_tiehi
XFILLER_37_216 VPWR VGND sg13g2_fill_1
XFILLER_19_975 VPWR VGND sg13g2_decap_8
X_4840_ _1689_ net1261 net392 VPWR VGND sg13g2_xnor2_1
X_4771_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[8\] _1630_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[9\]
+ _1631_ VPWR VGND sg13g2_nand3_1
X_6510_ net212 VGND VPWR net1362 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[11\]
+ clknet_leaf_44_clk sg13g2_dfrbpq_2
X_3722_ net404 _0685_ _0636_ _0775_ VPWR VGND sg13g2_nand3_1
X_6441_ net306 VGND VPWR net777 u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[7\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_1
X_3653_ _0706_ net406 _0660_ VPWR VGND sg13g2_xnor2_1
X_6372_ VGND VPWR net854 _2921_ _2924_ net916 sg13g2_a21oi_1
X_5323_ _2075_ VPWR _2078_ VGND _2071_ _2076_ sg13g2_o21ai_1
X_3584_ net546 u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[1\] u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[1\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[1\] net535 net544 _0637_
+ VPWR VGND sg13g2_mux4_1
X_5254_ _2024_ _2025_ _2023_ _2026_ VPWR VGND sg13g2_nand3_1
X_5185_ _1966_ net1062 _1964_ VPWR VGND sg13g2_xnor2_1
X_4205_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[1\] net382
+ _1160_ VPWR VGND sg13g2_nor2_1
X_4136_ _1102_ _1097_ _1099_ _1101_ VPWR VGND sg13g2_and3_1
X_4067_ net879 _0987_ _1053_ VPWR VGND sg13g2_nor2b_1
XFILLER_19_1017 VPWR VGND sg13g2_decap_8
XFILLER_24_444 VPWR VGND sg13g2_fill_2
XFILLER_25_945 VPWR VGND sg13g2_fill_1
XFILLER_19_1028 VPWR VGND sg13g2_fill_1
XFILLER_25_989 VPWR VGND sg13g2_decap_8
X_4969_ net467 VPWR _1797_ VGND _1794_ _1795_ sg13g2_o21ai_1
X_6708_ net717 VGND VPWR _0317_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[5\]\[4\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_1
X_6639_ net83 VGND VPWR _0248_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt_sum\[5\]
+ clknet_leaf_5_clk sg13g2_dfrbpq_2
Xheichips25_CORDIC_39 VPWR VGND uo_out[6] sg13g2_tielo
Xheichips25_CORDIC_28 VPWR VGND uio_oe[4] sg13g2_tielo
XFILLER_47_42 VPWR VGND sg13g2_fill_2
XFILLER_47_75 VPWR VGND sg13g2_decap_4
XFILLER_34_219 VPWR VGND sg13g2_fill_1
XFILLER_16_956 VPWR VGND sg13g2_decap_8
XFILLER_42_274 VPWR VGND sg13g2_fill_1
XFILLER_8_47 VPWR VGND sg13g2_fill_2
XFILLER_7_621 VPWR VGND sg13g2_fill_2
XFILLER_3_871 VPWR VGND sg13g2_decap_8
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk VPWR VGND sg13g2_buf_8
X_5941_ VGND VPWR _2596_ _2600_ _0396_ _2601_ sg13g2_a21oi_1
XFILLER_46_591 VPWR VGND sg13g2_fill_1
X_5872_ _2543_ net1422 _2541_ VPWR VGND sg13g2_xnor2_1
X_6577__145 VPWR VGND net145 sg13g2_tiehi
XFILLER_22_937 VPWR VGND sg13g2_decap_8
X_4823_ _1675_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[7\] net391
+ VPWR VGND sg13g2_xnor2_1
X_4754_ _1617_ net401 _1499_ VPWR VGND sg13g2_nand2b_1
X_3705_ _0756_ _0689_ _0758_ VPWR VGND sg13g2_xor2_1
X_4685_ net394 _1558_ _1559_ VPWR VGND sg13g2_and2_1
X_6424_ net332 VGND VPWR net921 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[2\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_2
X_3636_ _0689_ net406 _0688_ VPWR VGND sg13g2_nand2_1
X_3567_ u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[5\] u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[4\]
+ u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[6\] _0626_ VPWR VGND sg13g2_nand3_1
X_6669__53 VPWR VGND net53 sg13g2_tiehi
X_6355_ _2913_ net847 net880 _2910_ VPWR VGND sg13g2_and3_1
X_6286_ _2884_ _2883_ net402 VPWR VGND sg13g2_nand2b_1
XFILLER_1_819 VPWR VGND sg13g2_decap_8
X_5306_ net435 _2064_ net1269 _0297_ VPWR VGND sg13g2_nor3_1
X_3498_ _0568_ net1410 VPWR VGND sg13g2_inv_2
X_5237_ _2005_ _2011_ _2012_ VPWR VGND sg13g2_nor2b_1
XFILLER_25_1010 VPWR VGND sg13g2_decap_8
X_6584__138 VPWR VGND net138 sg13g2_tiehi
X_6746__495 VPWR VGND net679 sg13g2_tiehi
X_5168_ _1952_ net1291 net380 VPWR VGND sg13g2_xnor2_1
X_5099_ VGND VPWR net415 _1891_ _1892_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[2\]
+ sg13g2_a21oi_1
X_4119_ net1060 net533 _1088_ VPWR VGND sg13g2_xor2_1
XFILLER_13_937 VPWR VGND sg13g2_decap_8
XFILLER_24_285 VPWR VGND sg13g2_fill_1
XFILLER_12_469 VPWR VGND sg13g2_fill_1
X_6753__488 VPWR VGND net672 sg13g2_tiehi
XFILLER_3_112 VPWR VGND sg13g2_fill_1
XFILLER_0_885 VPWR VGND sg13g2_decap_8
Xhold7 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[2\] VPWR VGND net764
+ sg13g2_dlygate4sd3_1
XFILLER_28_591 VPWR VGND sg13g2_fill_1
XFILLER_8_930 VPWR VGND sg13g2_decap_8
XFILLER_12_970 VPWR VGND sg13g2_decap_8
XFILLER_31_789 VPWR VGND sg13g2_fill_1
XFILLER_7_462 VPWR VGND sg13g2_fill_1
Xhold407 _0268_ VPWR VGND net1164 sg13g2_dlygate4sd3_1
Xhold418 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[7\] VPWR VGND net1175
+ sg13g2_dlygate4sd3_1
X_4470_ _1380_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[1\]
+ _1379_ VPWR VGND sg13g2_xnor2_1
XFILLER_7_495 VPWR VGND sg13g2_fill_2
Xhold429 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[9\] VPWR VGND net1186
+ sg13g2_dlygate4sd3_1
XFILLER_48_1021 VPWR VGND sg13g2_decap_8
X_6140_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[5\] net416 _2758_
+ _2765_ VPWR VGND sg13g2_a21o_1
X_6071_ _2698_ VPWR _2706_ VGND net511 _0622_ sg13g2_o21ai_1
X_6666__56 VPWR VGND net56 sg13g2_tiehi
X_5022_ net1489 _1840_ _0238_ VPWR VGND sg13g2_nor2b_1
XFILLER_17_0 VPWR VGND sg13g2_fill_1
X_5924_ VPWR _2587_ _2586_ VGND sg13g2_inv_1
X_5855_ _0580_ _2527_ _2528_ VPWR VGND sg13g2_nor2_1
X_4806_ _1661_ net1237 net391 VPWR VGND sg13g2_nand2_1
XFILLER_9_90 VPWR VGND sg13g2_fill_1
XFILLER_10_929 VPWR VGND sg13g2_decap_8
X_5786_ _2465_ _2463_ _2461_ _2469_ VPWR VGND sg13g2_a21o_1
X_4737_ _1603_ net1458 net400 VPWR VGND sg13g2_nand2_1
X_4668_ _1545_ net1188 net394 VPWR VGND sg13g2_xnor2_1
X_6407_ net366 VGND VPWR net945 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[4\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
X_3619_ _0672_ _0640_ _0671_ VPWR VGND sg13g2_nand2_1
X_4599_ _1480_ VPWR _1487_ VGND _1482_ _1484_ sg13g2_o21ai_1
X_6338_ net374 _2901_ net932 _0504_ VPWR VGND sg13g2_nor3_1
X_6269_ net1070 VPWR _2870_ VGND _0543_ net939 sg13g2_o21ai_1
XFILLER_17_517 VPWR VGND sg13g2_fill_1
XFILLER_5_933 VPWR VGND sg13g2_decap_8
XFILLER_0_682 VPWR VGND sg13g2_decap_8
X_6567__155 VPWR VGND net155 sg13g2_tiehi
XFILLER_39_108 VPWR VGND sg13g2_fill_1
XFILLER_39_119 VPWR VGND sg13g2_fill_1
X_6663__59 VPWR VGND net59 sg13g2_tiehi
XFILLER_48_697 VPWR VGND sg13g2_fill_2
XFILLER_35_303 VPWR VGND sg13g2_fill_1
XFILLER_36_815 VPWR VGND sg13g2_fill_2
X_3970_ _0971_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[8\] _0964_
+ VPWR VGND sg13g2_xnor2_1
X_5640_ _2336_ net1258 _2347_ VPWR VGND sg13g2_xor2_1
X_6574__148 VPWR VGND net148 sg13g2_tiehi
X_5571_ _2285_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[3\]
+ _2287_ VPWR VGND sg13g2_xor2_1
XFILLER_31_597 VPWR VGND sg13g2_fill_2
X_4522_ net384 net1477 _1425_ VPWR VGND sg13g2_xor2_1
Xhold204 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[5\] VPWR VGND
+ net961 sg13g2_dlygate4sd3_1
Xhold226 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[10\] VPWR VGND net983 sg13g2_dlygate4sd3_1
XFILLER_8_793 VPWR VGND sg13g2_fill_2
Xhold215 _0300_ VPWR VGND net972 sg13g2_dlygate4sd3_1
X_4453_ _1367_ net486 _1366_ VPWR VGND sg13g2_nand2b_1
Xhold259 _0376_ VPWR VGND net1016 sg13g2_dlygate4sd3_1
Xhold248 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[2\] VPWR VGND net1005
+ sg13g2_dlygate4sd3_1
Xhold237 _1563_ VPWR VGND net994 sg13g2_dlygate4sd3_1
X_4384_ _1307_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[8\] _1306_
+ VPWR VGND sg13g2_xnor2_1
X_6123_ _2749_ _2750_ _0429_ VPWR VGND sg13g2_nor2b_1
X_6054_ net1522 _2690_ _2691_ VPWR VGND sg13g2_and2_1
X_5005_ net469 VPWR _1826_ VGND net988 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].y_shr\[0\]
+ sg13g2_o21ai_1
X_6743__498 VPWR VGND net682 sg13g2_tiehi
XFILLER_38_185 VPWR VGND sg13g2_fill_2
XFILLER_41_306 VPWR VGND sg13g2_fill_2
X_5907_ _2570_ net1509 _2572_ VPWR VGND sg13g2_xor2_1
X_6887_ net298 VGND VPWR net797 u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[7\]
+ clknet_leaf_13_clk sg13g2_dfrbpq_1
X_5838_ VGND VPWR _0577_ _2497_ _2513_ net514 sg13g2_a21oi_1
X_5769_ VGND VPWR net519 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[6\]
+ _2455_ _2453_ sg13g2_a21oi_1
XFILLER_2_914 VPWR VGND sg13g2_decap_8
Xhold760 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[2\] VPWR VGND net1517
+ sg13g2_dlygate4sd3_1
Xhold782 _2012_ VPWR VGND net1539 sg13g2_dlygate4sd3_1
Xhold771 _1250_ VPWR VGND net1528 sg13g2_dlygate4sd3_1
Xhold793 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[5\] VPWR VGND net1550
+ sg13g2_dlygate4sd3_1
XFILLER_9_535 VPWR VGND sg13g2_fill_2
X_6458__277 VPWR VGND net277 sg13g2_tiehi
XFILLER_5_730 VPWR VGND sg13g2_decap_8
XFILLER_4_284 VPWR VGND sg13g2_fill_1
XFILLER_1_980 VPWR VGND sg13g2_decap_8
X_6810_ net615 VGND VPWR net1211 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[5\]
+ clknet_leaf_63_clk sg13g2_dfrbpq_1
XFILLER_24_829 VPWR VGND sg13g2_fill_2
XFILLER_17_870 VPWR VGND sg13g2_fill_2
XFILLER_23_317 VPWR VGND sg13g2_fill_2
XFILLER_36_689 VPWR VGND sg13g2_fill_1
X_6741_ net684 VGND VPWR _0350_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[12\]
+ clknet_leaf_57_clk sg13g2_dfrbpq_2
X_3953_ _0954_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[14\] _0953_
+ VPWR VGND sg13g2_xnor2_1
X_3884_ _0908_ _0536_ _0904_ VPWR VGND sg13g2_xnor2_1
X_6672_ net50 VGND VPWR _0281_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[0\]
+ clknet_leaf_46_clk sg13g2_dfrbpq_2
X_5623_ net474 VPWR _2333_ VGND _2328_ _2332_ sg13g2_o21ai_1
X_5554_ _0593_ _2271_ _2272_ VPWR VGND sg13g2_nor2_1
X_5485_ _2218_ _0559_ _2206_ VPWR VGND sg13g2_xnor2_1
X_4505_ _1411_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[10\]
+ _1410_ VPWR VGND sg13g2_xnor2_1
X_4436_ VGND VPWR _1348_ _1351_ _0140_ _1352_ sg13g2_a21oi_1
Xfanout514 net1247 net514 VPWR VGND sg13g2_buf_8
X_4367_ _1295_ net503 _1294_ VPWR VGND sg13g2_nand2_1
Xfanout503 net504 net503 VPWR VGND sg13g2_buf_2
X_6106_ _2736_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[0\] net965
+ VPWR VGND sg13g2_xnor2_1
Xfanout525 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].z_sign net525
+ VPWR VGND sg13g2_buf_8
Xfanout547 u_angle_cordic_12b_pmod.waveform_sel_reg\[0\] net547 VPWR VGND sg13g2_buf_8
Xfanout536 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].z_sign net536
+ VPWR VGND sg13g2_buf_8
X_4298_ _1239_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[8\] net381
+ VPWR VGND sg13g2_xnor2_1
X_6037_ _2671_ VPWR _2676_ VGND _2667_ _2672_ sg13g2_o21ai_1
X_6557__165 VPWR VGND net165 sg13g2_tiehi
XFILLER_2_711 VPWR VGND sg13g2_decap_8
Xhold590 _2523_ VPWR VGND net1347 sg13g2_dlygate4sd3_1
XFILLER_2_788 VPWR VGND sg13g2_decap_8
X_6564__158 VPWR VGND net158 sg13g2_tiehi
XFILLER_12_1012 VPWR VGND sg13g2_decap_8
X_5270_ net528 net862 _2036_ VPWR VGND sg13g2_nor2b_1
X_4221_ _1165_ _1166_ _1169_ _1173_ VPWR VGND sg13g2_or3_1
X_4152_ _0094_ net504 _1113_ net1037 VPWR VGND sg13g2_and3_1
X_4083_ _0986_ _1062_ net824 _1064_ VPWR VGND sg13g2_nand3_1
X_4985_ _1810_ _1799_ _1808_ _1809_ VPWR VGND sg13g2_and3_1
X_6724_ net701 VGND VPWR net1157 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[7\]
+ clknet_leaf_30_clk sg13g2_dfrbpq_2
X_3936_ _0532_ net982 net1012 net918 _0938_ VPWR VGND sg13g2_nor4_1
X_3867_ _0895_ _0885_ _0894_ VPWR VGND sg13g2_nand2_1
X_6655_ net67 VGND VPWR net1395 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[2\]
+ clknet_leaf_48_clk sg13g2_dfrbpq_1
X_6586_ net136 VGND VPWR net1274 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[11\]
+ clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3798_ _0829_ _0842_ _0844_ _0845_ VPWR VGND sg13g2_nor3_1
X_5606_ VPWR _2318_ net1402 VGND sg13g2_inv_1
XFILLER_3_508 VPWR VGND sg13g2_fill_2
X_5537_ _2257_ _2258_ _2260_ VPWR VGND sg13g2_nor2_1
X_5468_ _2204_ _2203_ _2199_ VPWR VGND sg13g2_nand2b_1
X_5399_ net478 VPWR _2145_ VGND _2141_ _2144_ sg13g2_o21ai_1
X_4419_ _1338_ net1411 _1337_ VPWR VGND sg13g2_nand2_1
Xfanout388 net390 net388 VPWR VGND sg13g2_buf_8
Xfanout399 _1783_ net399 VPWR VGND sg13g2_buf_8
Xfanout377 net378 net377 VPWR VGND sg13g2_buf_8
XFILLER_36_33 VPWR VGND sg13g2_fill_2
XFILLER_36_55 VPWR VGND sg13g2_fill_1
XFILLER_43_946 VPWR VGND sg13g2_fill_1
XFILLER_11_898 VPWR VGND sg13g2_decap_8
XFILLER_7_869 VPWR VGND sg13g2_decap_8
XFILLER_42_1027 VPWR VGND sg13g2_fill_2
XFILLER_18_442 VPWR VGND sg13g2_fill_1
XFILLER_19_954 VPWR VGND sg13g2_decap_8
XFILLER_45_250 VPWR VGND sg13g2_fill_1
X_4770_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[7\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[6\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[5\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[9\]\[4\]
+ _1630_ VPWR VGND sg13g2_and4_1
XFILLER_14_692 VPWR VGND sg13g2_fill_1
XFILLER_9_140 VPWR VGND sg13g2_fill_2
X_3721_ VGND VPWR _0752_ _0758_ _0774_ _0757_ sg13g2_a21oi_1
X_6440_ net307 VGND VPWR net782 u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[6\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_1
X_3652_ VPWR _0705_ _0704_ VGND sg13g2_inv_1
X_6371_ VGND VPWR net854 _2921_ _0516_ _2923_ sg13g2_a21oi_1
X_3583_ u_angle_cordic_12b_pmod.waveform_sel_reg\[0\] u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[11\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[11\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[11\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp\[11\] net1514 _0636_
+ VPWR VGND sg13g2_mux4_1
X_5322_ VGND VPWR _2071_ _2076_ _0301_ _2077_ sg13g2_a21oi_1
X_5253_ _2007_ VPWR _2025_ VGND net1181 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[4\]
+ sg13g2_o21ai_1
X_5184_ _1965_ net1062 _1964_ VPWR VGND sg13g2_nand2_1
X_4204_ VGND VPWR net531 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[12\]
+ _1159_ _1153_ sg13g2_a21oi_1
X_4135_ net1149 net534 _1101_ VPWR VGND sg13g2_xor2_1
X_6547__175 VPWR VGND net175 sg13g2_tiehi
XFILLER_28_228 VPWR VGND sg13g2_fill_1
X_4066_ net449 net16 _0069_ VPWR VGND sg13g2_and2_1
XFILLER_25_968 VPWR VGND sg13g2_decap_8
XFILLER_24_489 VPWR VGND sg13g2_fill_1
X_4968_ VPWR _1796_ _1795_ VGND sg13g2_inv_1
X_4899_ net390 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[7\] _1738_
+ VPWR VGND sg13g2_xor2_1
X_3919_ net450 net781 _0049_ VPWR VGND sg13g2_and2_1
X_6707_ net718 VGND VPWR net1368 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[5\]\[3\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_1
X_6638_ net84 VGND VPWR net1198 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[11\]
+ clknet_leaf_24_clk sg13g2_dfrbpq_1
X_6554__168 VPWR VGND net168 sg13g2_tiehi
XFILLER_4_839 VPWR VGND sg13g2_decap_8
Xheichips25_CORDIC_29 VPWR VGND uio_oe[5] sg13g2_tielo
X_6569_ net153 VGND VPWR net1191 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[7\]
+ clknet_leaf_31_clk sg13g2_dfrbpq_2
XFILLER_47_537 VPWR VGND sg13g2_fill_2
XFILLER_47_54 VPWR VGND sg13g2_decap_8
XFILLER_19_217 VPWR VGND sg13g2_fill_1
XFILLER_16_935 VPWR VGND sg13g2_decap_8
XFILLER_43_721 VPWR VGND sg13g2_fill_1
X_6461__273 VPWR VGND net273 sg13g2_tiehi
X_6693__562 VPWR VGND net746 sg13g2_tiehi
XFILLER_7_611 VPWR VGND sg13g2_fill_2
XFILLER_3_850 VPWR VGND sg13g2_decap_8
X_5940_ net458 VPWR _2601_ VGND _2596_ _2600_ sg13g2_o21ai_1
X_5871_ _2542_ net1422 _2541_ VPWR VGND sg13g2_nand2_1
XFILLER_15_990 VPWR VGND sg13g2_decap_8
XFILLER_33_275 VPWR VGND sg13g2_fill_1
X_4822_ VGND VPWR net1091 net391 _1674_ _1672_ sg13g2_a21oi_1
X_4753_ _1616_ _1610_ _1613_ VPWR VGND sg13g2_nand2_1
X_3704_ _0689_ _0756_ _0757_ VPWR VGND sg13g2_nor2_1
X_6915__268 VPWR VGND net268 sg13g2_tiehi
X_6423_ net334 VGND VPWR net1025 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[1\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_2
X_4684_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[0\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[1\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[2\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[3\]
+ _1558_ VPWR VGND sg13g2_nor4_1
X_3635_ _0685_ net405 _0688_ VPWR VGND sg13g2_xor2_1
X_3566_ net878 net442 _0520_ VPWR VGND sg13g2_and2_1
X_6354_ VGND VPWR net847 _2910_ _0510_ _2912_ sg13g2_a21oi_1
X_6285_ _2883_ net1043 _2881_ VPWR VGND sg13g2_xnor2_1
X_3497_ _0567_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[10\]
+ VPWR VGND sg13g2_inv_2
X_5305_ VGND VPWR _2059_ _2061_ _2065_ _2063_ sg13g2_a21oi_1
X_5236_ _2011_ net1551 _2009_ VPWR VGND sg13g2_xnor2_1
X_5167_ _0272_ net493 _1950_ _1951_ VPWR VGND sg13g2_and3_1
X_5098_ VGND VPWR _1891_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[1\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[0\] sg13g2_or2_1
X_4118_ _1087_ _0582_ net1060 VPWR VGND sg13g2_nand2_1
XFILLER_44_529 VPWR VGND sg13g2_fill_2
X_4049_ _1040_ _1038_ _1041_ VPWR VGND sg13g2_nor2b_1
XFILLER_13_916 VPWR VGND sg13g2_decap_8
XFILLER_40_746 VPWR VGND sg13g2_fill_1
XFILLER_21_982 VPWR VGND sg13g2_decap_8
XFILLER_32_1026 VPWR VGND sg13g2_fill_2
XFILLER_20_492 VPWR VGND sg13g2_fill_1
XFILLER_0_864 VPWR VGND sg13g2_decap_8
Xhold8 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[0\]\[0\] VPWR VGND net765
+ sg13g2_dlygate4sd3_1
XFILLER_30_289 VPWR VGND sg13g2_fill_2
Xhold408 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[1\] VPWR VGND net1165
+ sg13g2_dlygate4sd3_1
XFILLER_8_986 VPWR VGND sg13g2_decap_8
X_6537__185 VPWR VGND net185 sg13g2_tiehi
Xhold419 _0090_ VPWR VGND net1176 sg13g2_dlygate4sd3_1
X_6070_ _2703_ _2705_ _0421_ VPWR VGND sg13g2_nor2_1
X_5021_ VGND VPWR _1832_ _1838_ _1840_ net427 sg13g2_a21oi_1
XFILLER_39_824 VPWR VGND sg13g2_fill_2
XFILLER_26_518 VPWR VGND sg13g2_fill_2
XFILLER_38_367 VPWR VGND sg13g2_fill_1
X_6544__178 VPWR VGND net178 sg13g2_tiehi
X_5923_ _2586_ net1381 _2584_ VPWR VGND sg13g2_xnor2_1
X_5854_ _2527_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[8\]
+ _2526_ VPWR VGND sg13g2_xnor2_1
X_4805_ VGND VPWR _1653_ _1660_ net1569 net536 sg13g2_a21oi_2
XFILLER_10_908 VPWR VGND sg13g2_decap_8
X_5785_ _2467_ _2468_ _0373_ VPWR VGND sg13g2_nor2_1
X_4736_ _1596_ _1600_ _1602_ VPWR VGND sg13g2_nor2_1
X_6590__132 VPWR VGND net132 sg13g2_tiehi
X_4667_ VGND VPWR net1017 net393 _1544_ _1543_ sg13g2_a21oi_1
X_6406_ net368 VGND VPWR net911 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[3\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
X_3618_ net403 net405 _0671_ VPWR VGND sg13g2_xor2_1
X_4598_ net437 _1485_ _1486_ _0168_ VPWR VGND sg13g2_nor3_1
X_6337_ net931 _2899_ _2902_ VPWR VGND sg13g2_nor2_1
XFILLER_0_105 VPWR VGND sg13g2_fill_1
X_3549_ VPWR _0619_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[3\] VGND
+ sg13g2_inv_1
X_6268_ _2868_ _2869_ _2866_ _0458_ VPWR VGND sg13g2_mux2_1
X_5219_ net439 _1995_ _0280_ VPWR VGND sg13g2_nor2_1
X_6199_ _2816_ net1281 _2817_ VPWR VGND sg13g2_xor2_1
X_6683__572 VPWR VGND net756 sg13g2_tiehi
XFILLER_13_702 VPWR VGND sg13g2_fill_2
XFILLER_8_205 VPWR VGND sg13g2_fill_1
XFILLER_5_912 VPWR VGND sg13g2_decap_8
X_6690__565 VPWR VGND net749 sg13g2_tiehi
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk VPWR VGND sg13g2_buf_8
XFILLER_5_989 VPWR VGND sg13g2_decap_8
XFILLER_0_661 VPWR VGND sg13g2_decap_8
X_5570_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[3\] _2285_
+ _2286_ VPWR VGND sg13g2_nor2_1
X_4521_ VGND VPWR _1421_ _1423_ _0153_ _1424_ sg13g2_a21oi_1
XFILLER_7_293 VPWR VGND sg13g2_fill_1
XFILLER_7_282 VPWR VGND sg13g2_fill_1
Xhold216 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[2\]\[0\] VPWR VGND net973
+ sg13g2_dlygate4sd3_1
Xhold205 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[0\] VPWR VGND net962
+ sg13g2_dlygate4sd3_1
X_4452_ _1365_ _1364_ _1366_ VPWR VGND sg13g2_nor2b_1
Xhold249 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[1\] VPWR VGND net1006
+ sg13g2_dlygate4sd3_1
Xhold227 _0030_ VPWR VGND net984 sg13g2_dlygate4sd3_1
Xhold238 _0184_ VPWR VGND net995 sg13g2_dlygate4sd3_1
X_4383_ net542 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[7\] _1306_
+ VPWR VGND sg13g2_nor2b_1
X_6122_ VGND VPWR _2742_ _2748_ _2750_ net422 sg13g2_a21oi_1
X_6053_ _2690_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[6\]
+ _2689_ VPWR VGND sg13g2_xnor2_1
X_5004_ _1825_ net988 net1052 VPWR VGND sg13g2_nand2_1
XFILLER_22_1014 VPWR VGND sg13g2_decap_8
X_6662__60 VPWR VGND net60 sg13g2_tiehi
X_5906_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[1\] _2570_
+ _2571_ VPWR VGND sg13g2_and2_1
XFILLER_22_510 VPWR VGND sg13g2_fill_2
X_6886_ net300 VGND VPWR _0495_ u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[6\]
+ clknet_leaf_27_clk sg13g2_dfrbpq_1
X_5837_ _2507_ _2503_ _2506_ _2512_ VPWR VGND sg13g2_a21o_1
XFILLER_6_709 VPWR VGND sg13g2_decap_8
X_5768_ _2453_ _2454_ _0370_ VPWR VGND sg13g2_nor2b_1
X_4719_ _1588_ net1524 _1585_ VPWR VGND sg13g2_xnor2_1
X_5699_ VPWR _2398_ _2397_ VGND sg13g2_inv_1
Xhold761 _0302_ VPWR VGND net1518 sg13g2_dlygate4sd3_1
Xhold772 _0118_ VPWR VGND net1529 sg13g2_dlygate4sd3_1
Xhold750 _2256_ VPWR VGND net1507 sg13g2_dlygate4sd3_1
Xhold794 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[2\] VPWR
+ VGND net1551 sg13g2_dlygate4sd3_1
Xhold783 _0282_ VPWR VGND net1540 sg13g2_dlygate4sd3_1
X_6527__195 VPWR VGND net195 sg13g2_tiehi
X_6534__188 VPWR VGND net188 sg13g2_tiehi
XFILLER_5_786 VPWR VGND sg13g2_decap_8
XFILLER_48_451 VPWR VGND sg13g2_fill_1
XFILLER_48_484 VPWR VGND sg13g2_fill_1
X_6580__142 VPWR VGND net142 sg13g2_tiehi
XFILLER_24_819 VPWR VGND sg13g2_fill_2
X_6740_ net685 VGND VPWR net1195 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[11\]
+ clknet_leaf_57_clk sg13g2_dfrbpq_2
X_3952_ _0947_ _0952_ _0953_ VPWR VGND sg13g2_nor2b_1
X_3883_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[1\] u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[0\]
+ net920 _0907_ VPWR VGND sg13g2_nand3_1
X_6671_ net51 VGND VPWR _0280_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[6\]\[5\]
+ clknet_leaf_51_clk sg13g2_dfrbpq_1
XFILLER_31_351 VPWR VGND sg13g2_fill_2
X_5622_ _2332_ _0599_ _2330_ VPWR VGND sg13g2_xnor2_1
X_5553_ _2271_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[1\]
+ _2270_ VPWR VGND sg13g2_xnor2_1
X_4504_ net543 _1403_ _1410_ VPWR VGND sg13g2_nor2_1
X_5484_ _0323_ net479 _2216_ _2217_ VPWR VGND sg13g2_and3_1
X_4435_ net487 VPWR _1352_ VGND _1348_ _1351_ sg13g2_o21ai_1
Xfanout515 net516 net515 VPWR VGND sg13g2_buf_8
Xfanout504 net505 net504 VPWR VGND sg13g2_buf_8
X_4366_ VGND VPWR _1294_ _1293_ _1292_ sg13g2_or2_1
Xfanout537 net538 net537 VPWR VGND sg13g2_buf_2
X_6105_ net1046 _0545_ _2735_ VPWR VGND sg13g2_nor2_1
Xfanout526 net530 net526 VPWR VGND sg13g2_buf_8
Xfanout548 net551 net548 VPWR VGND sg13g2_buf_2
X_4297_ net437 net1463 _1238_ _0115_ VPWR VGND sg13g2_nor3_1
X_6036_ _2671_ _2673_ _2675_ VPWR VGND sg13g2_and2_1
XFILLER_26_145 VPWR VGND sg13g2_fill_1
X_6869_ net347 VGND VPWR _0478_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[1\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_2_767 VPWR VGND sg13g2_decap_8
XFILLER_1_222 VPWR VGND sg13g2_fill_1
Xhold580 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[5\]\[2\] VPWR VGND net1337
+ sg13g2_dlygate4sd3_1
Xhold591 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[4\] VPWR VGND net1348
+ sg13g2_dlygate4sd3_1
XFILLER_14_885 VPWR VGND sg13g2_decap_8
XFILLER_40_181 VPWR VGND sg13g2_fill_1
XFILLER_9_399 VPWR VGND sg13g2_fill_2
X_6395__387 VPWR VGND net571 sg13g2_tiehi
X_6471__253 VPWR VGND net253 sg13g2_tiehi
X_4220_ _1172_ net1300 net383 VPWR VGND sg13g2_xnor2_1
X_4151_ _0582_ VPWR _1114_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[9\]
+ net1036 sg13g2_o21ai_1
X_4082_ _1062_ _0987_ net824 _1063_ VPWR VGND sg13g2_a21o_1
XFILLER_48_292 VPWR VGND sg13g2_fill_1
X_4984_ net397 VPWR _1809_ VGND net1122 net1433 sg13g2_o21ai_1
XFILLER_23_148 VPWR VGND sg13g2_fill_2
X_6723_ net702 VGND VPWR _0332_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[6\]
+ clknet_leaf_30_clk sg13g2_dfrbpq_2
X_3935_ _0937_ net885 net548 VPWR VGND sg13g2_nand2b_1
X_6654_ net68 VGND VPWR net1102 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[1\]
+ clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_32_682 VPWR VGND sg13g2_fill_1
X_3866_ net842 _0890_ net887 _0894_ VPWR VGND sg13g2_nand3_1
X_5605_ _2317_ net1401 _2315_ VPWR VGND sg13g2_xnor2_1
X_6585_ net137 VGND VPWR _0194_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[10\]
+ clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3797_ _0832_ _0833_ _0831_ _0844_ VPWR VGND _0843_ sg13g2_nand4_1
X_5536_ _2257_ _2258_ _2259_ VPWR VGND sg13g2_and2_1
X_5467_ _2203_ net1502 _2201_ VPWR VGND sg13g2_xnor2_1
X_4418_ _1335_ _1336_ _1337_ VPWR VGND sg13g2_nor2b_1
X_5398_ _2144_ _2143_ _2142_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_1020 VPWR VGND sg13g2_decap_8
X_4349_ net436 _1278_ _1279_ _0126_ VPWR VGND sg13g2_nor3_1
Xfanout389 net390 net389 VPWR VGND sg13g2_buf_8
Xfanout378 _0988_ net378 VPWR VGND sg13g2_buf_2
X_6019_ net416 VPWR _2660_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[0\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[1\] sg13g2_o21ai_1
XFILLER_15_627 VPWR VGND sg13g2_fill_2
XFILLER_28_999 VPWR VGND sg13g2_decap_8
X_6524__198 VPWR VGND net198 sg13g2_tiehi
XFILLER_14_159 VPWR VGND sg13g2_fill_2
XFILLER_7_848 VPWR VGND sg13g2_decap_8
XFILLER_11_877 VPWR VGND sg13g2_decap_8
X_6570__152 VPWR VGND net152 sg13g2_tiehi
XFILLER_7_0 VPWR VGND sg13g2_fill_2
XFILLER_19_933 VPWR VGND sg13g2_decap_8
XFILLER_18_487 VPWR VGND sg13g2_fill_2
XFILLER_42_991 VPWR VGND sg13g2_fill_2
XFILLER_20_118 VPWR VGND sg13g2_fill_2
X_3720_ _0773_ _0760_ _0762_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_40_clk clknet_4_15_0_clk clknet_leaf_40_clk VPWR VGND sg13g2_buf_8
X_3651_ _0704_ net406 _0660_ VPWR VGND sg13g2_nand2_1
X_6370_ net377 VPWR _2923_ VGND net854 _2921_ sg13g2_o21ai_1
X_3582_ net442 net822 _0634_ _0635_ _0003_ VPWR VGND sg13g2_and4_1
XFILLER_6_881 VPWR VGND sg13g2_decap_8
X_5321_ net477 VPWR _2077_ VGND _2071_ _2076_ sg13g2_o21ai_1
X_5252_ _2024_ _2019_ _2017_ VPWR VGND sg13g2_nand2b_1
X_6848__393 VPWR VGND net577 sg13g2_tiehi
X_5183_ _1964_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[6\] _1963_
+ VPWR VGND sg13g2_xnor2_1
X_4203_ VGND VPWR _1151_ _1156_ _0101_ _1158_ sg13g2_a21oi_1
X_4134_ VGND VPWR _1096_ _1098_ _0090_ _1100_ sg13g2_a21oi_1
XFILLER_3_1011 VPWR VGND sg13g2_decap_8
X_4065_ net449 net15 _0068_ VPWR VGND sg13g2_and2_1
XFILLER_33_991 VPWR VGND sg13g2_fill_1
X_4967_ _1795_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[5\] net397
+ VPWR VGND sg13g2_xnor2_1
X_4898_ _1737_ _1733_ _1735_ VPWR VGND sg13g2_nand2_1
X_3918_ net463 net808 _0048_ VPWR VGND sg13g2_and2_1
X_6706_ net719 VGND VPWR _0315_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[5\]\[2\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_1
XFILLER_20_641 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_31_clk clknet_4_9_0_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
X_6637_ net85 VGND VPWR _0246_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[10\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_1
X_3849_ net441 VPWR _0882_ VGND net1023 _0880_ sg13g2_o21ai_1
X_6568_ net154 VGND VPWR net1254 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[6\]
+ clknet_leaf_29_clk sg13g2_dfrbpq_2
XFILLER_4_818 VPWR VGND sg13g2_decap_8
X_5519_ net523 net1563 _2245_ VPWR VGND sg13g2_and2_1
X_6499_ net223 VGND VPWR net964 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[0\]
+ clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_16_914 VPWR VGND sg13g2_decap_8
XFILLER_28_774 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_22_clk clknet_4_7_0_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
XFILLER_7_623 VPWR VGND sg13g2_fill_1
X_6678__44 VPWR VGND net44 sg13g2_tiehi
XFILLER_38_527 VPWR VGND sg13g2_fill_2
X_5870_ _2541_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[10\]
+ _2540_ VPWR VGND sg13g2_xnor2_1
XFILLER_34_744 VPWR VGND sg13g2_fill_2
XFILLER_34_766 VPWR VGND sg13g2_fill_2
X_4821_ _1672_ _1673_ _0204_ VPWR VGND sg13g2_nor2_1
X_6891__542 VPWR VGND net726 sg13g2_tiehi
X_4752_ net400 net1273 _1615_ VPWR VGND sg13g2_xor2_1
Xclkbuf_leaf_13_clk clknet_4_6_0_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_3703_ _0756_ net407 _0754_ VPWR VGND sg13g2_xnor2_1
X_4683_ _1547_ _1548_ _1557_ VPWR VGND sg13g2_nor2_1
X_6422_ net336 VGND VPWR _0031_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[0\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_2
X_3634_ VGND VPWR _0687_ _0685_ net404 sg13g2_or2_1
X_3565_ net865 net444 _0530_ VPWR VGND sg13g2_and2_1
X_6353_ net378 VPWR _2912_ VGND net847 _2910_ sg13g2_o21ai_1
X_6284_ _2882_ net1043 _2881_ VPWR VGND sg13g2_nand2_2
X_3496_ VPWR _0566_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[5\]
+ VGND sg13g2_inv_1
X_5304_ _2064_ _2059_ _2061_ _2063_ VPWR VGND sg13g2_and3_1
X_5235_ net1551 _2009_ _2010_ VPWR VGND sg13g2_and2_1
X_5166_ _1949_ _1948_ _1947_ _1951_ VPWR VGND sg13g2_a21o_1
XFILLER_29_527 VPWR VGND sg13g2_decap_4
X_5097_ _1887_ VPWR _1890_ VGND _1883_ _1888_ sg13g2_o21ai_1
X_4117_ _1082_ _1085_ _1086_ VPWR VGND sg13g2_and2_1
XFILLER_44_508 VPWR VGND sg13g2_fill_1
X_4048_ _1040_ _1037_ _1039_ VPWR VGND sg13g2_nand2_1
X_6560__162 VPWR VGND net162 sg13g2_tiehi
X_5999_ VGND VPWR _2645_ _2644_ _2643_ sg13g2_or2_1
XFILLER_21_961 VPWR VGND sg13g2_decap_8
X_6675__47 VPWR VGND net47 sg13g2_tiehi
XFILLER_0_843 VPWR VGND sg13g2_decap_8
Xhold9 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[2\] VPWR VGND net766
+ sg13g2_dlygate4sd3_1
XFILLER_16_744 VPWR VGND sg13g2_fill_1
XFILLER_31_769 VPWR VGND sg13g2_fill_2
XFILLER_8_965 VPWR VGND sg13g2_decap_8
Xhold409 _0172_ VPWR VGND net1166 sg13g2_dlygate4sd3_1
X_5020_ _1832_ _1838_ _1839_ VPWR VGND sg13g2_nor2_1
XFILLER_31_4 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_2_clk clknet_4_1_0_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
X_6845__396 VPWR VGND net580 sg13g2_tiehi
XFILLER_0_1025 VPWR VGND sg13g2_decap_4
X_5922_ net1381 _2584_ _2585_ VPWR VGND sg13g2_and2_1
X_5853_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[7\] net413
+ _2520_ _2526_ VPWR VGND sg13g2_a21o_1
X_4804_ _0201_ net483 _1658_ _1659_ VPWR VGND sg13g2_and3_1
X_5784_ _2468_ net476 _2466_ VPWR VGND sg13g2_nand2_1
XFILLER_34_596 VPWR VGND sg13g2_fill_1
X_4735_ _1600_ _1601_ _0190_ VPWR VGND sg13g2_nor2_1
X_4666_ net432 _1542_ _1543_ _0179_ VPWR VGND sg13g2_nor3_1
X_6405_ net370 VGND VPWR net894 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[2\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
X_3617_ VPWR _0670_ _0669_ VGND sg13g2_inv_1
X_4597_ _1486_ _1480_ _1482_ _1484_ VPWR VGND sg13g2_and3_1
X_3548_ VPWR _0618_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[4\] VGND
+ sg13g2_inv_1
X_6336_ net931 _2899_ _2901_ VPWR VGND sg13g2_and2_1
X_3479_ VPWR _0549_ net909 VGND sg13g2_inv_1
X_6267_ net421 _2867_ _2869_ VPWR VGND sg13g2_nor2_1
X_5218_ _1995_ _1990_ _1994_ VPWR VGND sg13g2_xnor2_1
X_6198_ _2809_ net510 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[12\]
+ _2816_ VPWR VGND sg13g2_mux2_1
X_5149_ net1410 _1936_ _1937_ VPWR VGND sg13g2_and2_1
XFILLER_13_758 VPWR VGND sg13g2_fill_1
XFILLER_5_968 VPWR VGND sg13g2_decap_8
XFILLER_0_640 VPWR VGND sg13g2_fill_2
XFILLER_48_699 VPWR VGND sg13g2_fill_1
XFILLER_47_176 VPWR VGND sg13g2_fill_2
XFILLER_43_393 VPWR VGND sg13g2_fill_1
XFILLER_15_1011 VPWR VGND sg13g2_decap_8
XFILLER_31_599 VPWR VGND sg13g2_fill_1
X_4520_ net498 VPWR _1424_ VGND _1421_ _1423_ sg13g2_o21ai_1
XFILLER_8_795 VPWR VGND sg13g2_fill_1
Xhold217 _2555_ VPWR VGND net974 sg13g2_dlygate4sd3_1
Xhold206 _1188_ VPWR VGND net963 sg13g2_dlygate4sd3_1
X_4451_ _1365_ net1158 net386 VPWR VGND sg13g2_xnor2_1
Xhold228 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[0\] VPWR VGND net985
+ sg13g2_dlygate4sd3_1
Xhold239 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[0\] VPWR
+ VGND net996 sg13g2_dlygate4sd3_1
X_6550__172 VPWR VGND net172 sg13g2_tiehi
X_4382_ net435 net923 _0133_ VPWR VGND sg13g2_nor2_1
X_6121_ _2742_ _2748_ _2749_ VPWR VGND sg13g2_nor2_1
X_6052_ VGND VPWR net416 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[5\]
+ _2689_ _2684_ sg13g2_a21oi_1
XFILLER_22_0 VPWR VGND sg13g2_fill_2
X_5003_ VGND VPWR _1822_ _1823_ _0235_ _1824_ sg13g2_a21oi_1
XFILLER_27_806 VPWR VGND sg13g2_fill_2
XFILLER_38_187 VPWR VGND sg13g2_fill_1
X_5905_ _2570_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[5\] _2569_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_35_861 VPWR VGND sg13g2_fill_2
XFILLER_34_382 VPWR VGND sg13g2_fill_2
X_6885_ net315 VGND VPWR _0494_ u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[5\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_1
X_5836_ VGND VPWR _2503_ _2507_ _2511_ _2506_ sg13g2_a21oi_1
X_5767_ VGND VPWR _2451_ _2452_ _2454_ net427 sg13g2_a21oi_1
X_4718_ VPWR _1587_ _1586_ VGND sg13g2_inv_1
X_5698_ _2397_ _0595_ _2395_ VPWR VGND sg13g2_xnor2_1
X_4649_ _1520_ _1525_ _1529_ VPWR VGND sg13g2_nor2_1
XFILLER_30_69 VPWR VGND sg13g2_fill_1
XFILLER_2_949 VPWR VGND sg13g2_decap_8
Xhold740 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[8\] VPWR VGND net1497
+ sg13g2_dlygate4sd3_1
Xhold762 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[4\] VPWR
+ VGND net1519 sg13g2_dlygate4sd3_1
Xhold751 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[9\] VPWR
+ VGND net1508 sg13g2_dlygate4sd3_1
Xhold773 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[8\] VPWR
+ VGND net1530 sg13g2_dlygate4sd3_1
X_6319_ net465 net802 _0490_ VPWR VGND sg13g2_and2_1
Xhold784 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[6\] VPWR VGND net1541
+ sg13g2_dlygate4sd3_1
Xhold795 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[1\] VPWR
+ VGND net1552 sg13g2_dlygate4sd3_1
XFILLER_7_1009 VPWR VGND sg13g2_decap_8
XFILLER_44_135 VPWR VGND sg13g2_fill_2
XFILLER_13_544 VPWR VGND sg13g2_fill_1
XFILLER_25_371 VPWR VGND sg13g2_fill_2
XFILLER_5_765 VPWR VGND sg13g2_decap_8
X_6842__399 VPWR VGND net583 sg13g2_tiehi
XFILLER_23_319 VPWR VGND sg13g2_fill_1
X_3951_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[9\] VPWR _0952_
+ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[8\] _0946_ sg13g2_o21ai_1
X_6738__503 VPWR VGND net687 sg13g2_tiehi
X_6670_ net52 VGND VPWR _0279_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[6\]\[4\]
+ clknet_leaf_51_clk sg13g2_dfrbpq_1
X_3882_ _0906_ net920 _0885_ VPWR VGND sg13g2_nand2_1
X_5621_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[9\] _2330_ _2331_
+ VPWR VGND sg13g2_and2_1
X_5552_ net515 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[0\]
+ _2270_ VPWR VGND sg13g2_nor2b_1
X_4503_ VGND VPWR _1401_ _1406_ _1409_ _1405_ sg13g2_a21oi_1
X_5483_ _2215_ _2213_ _2212_ _2217_ VPWR VGND sg13g2_a21o_1
X_4434_ _1349_ _1350_ _1351_ VPWR VGND sg13g2_and2_1
Xfanout505 net851 net505 VPWR VGND sg13g2_buf_8
X_4365_ net1110 net541 _1293_ VPWR VGND sg13g2_xor2_1
X_6104_ VGND VPWR _2731_ _2733_ _0426_ _2734_ sg13g2_a21oi_1
Xfanout516 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].z_sign net516
+ VPWR VGND sg13g2_buf_8
Xfanout527 net530 net527 VPWR VGND sg13g2_buf_1
Xfanout538 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].z_sign net538
+ VPWR VGND sg13g2_buf_1
X_6035_ VGND VPWR _2667_ _2672_ _0417_ _2674_ sg13g2_a21oi_1
X_4296_ _1232_ _1236_ _1238_ VPWR VGND sg13g2_nor2b_1
Xfanout549 net551 net549 VPWR VGND sg13g2_buf_8
XFILLER_27_625 VPWR VGND sg13g2_fill_2
XFILLER_39_485 VPWR VGND sg13g2_fill_2
X_6868_ net349 VGND VPWR _0477_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[0\]
+ clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_34_190 VPWR VGND sg13g2_fill_2
X_5819_ net512 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[3\]
+ _2496_ VPWR VGND sg13g2_nor2b_1
X_6799_ net626 VGND VPWR _0408_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[6\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_2_746 VPWR VGND sg13g2_decap_8
Xhold570 _2537_ VPWR VGND net1327 sg13g2_dlygate4sd3_1
Xhold581 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[3\] VPWR VGND net1338
+ sg13g2_dlygate4sd3_1
Xhold592 _0380_ VPWR VGND net1349 sg13g2_dlygate4sd3_1
X_6865__355 VPWR VGND net355 sg13g2_tiehi
XFILLER_45_433 VPWR VGND sg13g2_fill_2
XFILLER_17_146 VPWR VGND sg13g2_fill_2
X_6540__182 VPWR VGND net182 sg13g2_tiehi
XFILLER_49_5 VPWR VGND sg13g2_decap_8
X_4150_ _1113_ _1111_ _1108_ VPWR VGND sg13g2_nand2b_1
XFILLER_49_750 VPWR VGND sg13g2_fill_2
X_4081_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[4\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[3\]
+ _1057_ _1062_ VPWR VGND sg13g2_or3_1
X_4983_ _1807_ VPWR _1808_ VGND net1433 net397 sg13g2_o21ai_1
X_3934_ VGND VPWR net961 _0935_ _0936_ net952 sg13g2_a21oi_1
X_6722_ net703 VGND VPWR net1359 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[5\]
+ clknet_leaf_47_clk sg13g2_dfrbpq_1
X_3865_ VGND VPWR net842 _0890_ _0893_ net887 sg13g2_a21oi_1
X_6653_ net69 VGND VPWR net1035 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[0\]
+ clknet_leaf_46_clk sg13g2_dfrbpq_1
X_5604_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[7\] _2315_ _2316_
+ VPWR VGND sg13g2_and2_1
X_6584_ net138 VGND VPWR _0193_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[9\]
+ clknet_leaf_34_clk sg13g2_dfrbpq_2
XFILLER_9_890 VPWR VGND sg13g2_decap_8
X_3796_ _0843_ _0551_ net1056 net892 _0536_ VPWR VGND sg13g2_a22oi_1
X_5535_ net1124 net523 _2258_ VPWR VGND sg13g2_xor2_1
X_5466_ _2202_ net1502 _2201_ VPWR VGND sg13g2_nand2_1
X_4417_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[12\] VPWR _1336_ VGND
+ net543 _1328_ sg13g2_o21ai_1
X_5397_ _2143_ net1386 _2132_ VPWR VGND sg13g2_nand2_1
X_4348_ _1279_ _1273_ _1275_ _1277_ VPWR VGND sg13g2_and3_1
Xfanout379 _2007_ net379 VPWR VGND sg13g2_buf_8
X_4279_ VGND VPWR _1217_ _1221_ _0113_ _1222_ sg13g2_a21oi_1
X_6018_ _2656_ VPWR _2659_ VGND _2652_ _2657_ sg13g2_o21ai_1
XFILLER_23_661 VPWR VGND sg13g2_fill_2
XFILLER_7_827 VPWR VGND sg13g2_decap_8
X_6728__513 VPWR VGND net697 sg13g2_tiehi
XFILLER_19_912 VPWR VGND sg13g2_decap_8
XFILLER_19_989 VPWR VGND sg13g2_decap_8
X_6735__506 VPWR VGND net690 sg13g2_tiehi
XFILLER_9_142 VPWR VGND sg13g2_fill_1
X_3650_ _0643_ net406 _0703_ VPWR VGND sg13g2_and2_1
X_3581_ VGND VPWR _0634_ net860 _0002_ _0633_ sg13g2_a21oi_1
XFILLER_6_860 VPWR VGND sg13g2_decap_8
X_5320_ _2076_ _0554_ _2074_ VPWR VGND sg13g2_xnor2_1
X_5251_ _2023_ net1227 net379 VPWR VGND sg13g2_xnor2_1
X_4202_ _1158_ net496 _1157_ VPWR VGND sg13g2_nand2_1
X_5182_ net526 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[5\] _1963_
+ VPWR VGND sg13g2_nor2b_1
XFILLER_3_83 VPWR VGND sg13g2_fill_2
X_4133_ _1100_ net501 _1099_ VPWR VGND sg13g2_nand2_1
X_4064_ _1051_ _1052_ _0067_ VPWR VGND sg13g2_nor2b_1
X_4966_ VGND VPWR net1112 net398 _1794_ _1792_ sg13g2_a21oi_1
X_6705_ net720 VGND VPWR net1305 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[5\]\[1\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_1
X_4897_ _1736_ _1735_ _0217_ VPWR VGND sg13g2_nor2b_1
X_3917_ net463 net805 _0047_ VPWR VGND sg13g2_and2_1
X_6855__376 VPWR VGND net560 sg13g2_tiehi
XFILLER_32_480 VPWR VGND sg13g2_fill_1
X_6636_ net86 VGND VPWR _0245_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[9\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_1
X_3848_ net1023 _0880_ _0881_ VPWR VGND sg13g2_and2_1
X_3779_ VGND VPWR _0540_ _0541_ _0827_ _0627_ sg13g2_a21oi_1
X_6567_ net155 VGND VPWR _0176_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[5\]
+ clknet_leaf_31_clk sg13g2_dfrbpq_1
X_5518_ net523 net1563 _2244_ VPWR VGND sg13g2_nor2_1
X_6498_ net224 VGND VPWR net1310 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[10\]
+ clknet_leaf_41_clk sg13g2_dfrbpq_2
X_5449_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[9\] net418 _2179_
+ _2187_ VPWR VGND sg13g2_a21o_1
X_6530__192 VPWR VGND net192 sg13g2_tiehi
XFILLER_47_23 VPWR VGND sg13g2_decap_8
XFILLER_42_211 VPWR VGND sg13g2_fill_1
XFILLER_24_981 VPWR VGND sg13g2_decap_8
XFILLER_10_130 VPWR VGND sg13g2_fill_2
XFILLER_6_123 VPWR VGND sg13g2_fill_1
XFILLER_3_885 VPWR VGND sg13g2_decap_8
XFILLER_33_8 VPWR VGND sg13g2_fill_1
XFILLER_33_233 VPWR VGND sg13g2_fill_2
X_4820_ net468 VPWR _1673_ VGND _1669_ _1671_ sg13g2_o21ai_1
X_4751_ VGND VPWR _1612_ _1613_ _0193_ _1614_ sg13g2_a21oi_1
X_3702_ VPWR _0755_ _0754_ VGND sg13g2_inv_1
X_4682_ VGND VPWR _1553_ _1555_ _0182_ _1556_ sg13g2_a21oi_1
X_6421_ net338 VGND VPWR net984 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[10\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
X_3633_ _0686_ net404 _0685_ VPWR VGND sg13g2_nand2_1
X_3564_ net821 net445 _0529_ VPWR VGND sg13g2_and2_1
X_6352_ net374 _2910_ net957 _0509_ VPWR VGND sg13g2_nor3_1
X_6283_ _2881_ net1041 net506 VPWR VGND sg13g2_nand2_2
X_3495_ _0565_ net1181 VPWR VGND sg13g2_inv_2
X_5303_ net1268 net529 _2063_ VPWR VGND sg13g2_xor2_1
X_5234_ net379 _2008_ _2009_ VPWR VGND sg13g2_and2_1
X_5165_ _1948_ _1949_ _1947_ _1950_ VPWR VGND sg13g2_nand3_1
XFILLER_25_1024 VPWR VGND sg13g2_decap_4
X_4116_ _0087_ net499 _1084_ _1085_ VPWR VGND sg13g2_and3_1
X_5096_ VGND VPWR _1883_ _1888_ _0263_ _1889_ sg13g2_a21oi_1
X_4047_ _1039_ net548 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[9\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_24_200 VPWR VGND sg13g2_fill_2
X_5998_ net1154 net513 _2644_ VPWR VGND sg13g2_xor2_1
X_4949_ _1780_ net1464 _1778_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_940 VPWR VGND sg13g2_decap_8
X_6718__523 VPWR VGND net707 sg13g2_tiehi
XFILLER_32_1028 VPWR VGND sg13g2_fill_1
X_6619_ net103 VGND VPWR _0228_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[4\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_0_822 VPWR VGND sg13g2_decap_8
XFILLER_0_899 VPWR VGND sg13g2_decap_8
X_6725__516 VPWR VGND net700 sg13g2_tiehi
XFILLER_8_944 VPWR VGND sg13g2_decap_8
X_6732__509 VPWR VGND net693 sg13g2_tiehi
XFILLER_12_984 VPWR VGND sg13g2_decap_8
X_6914__270 VPWR VGND net270 sg13g2_tiehi
XFILLER_3_682 VPWR VGND sg13g2_decap_8
XFILLER_2_192 VPWR VGND sg13g2_fill_2
X_6468__259 VPWR VGND net259 sg13g2_tiehi
X_5921_ _2584_ net1346 _2583_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_1004 VPWR VGND sg13g2_decap_8
XFILLER_46_380 VPWR VGND sg13g2_fill_1
X_5852_ _2522_ VPWR _2525_ VGND _2519_ _2523_ sg13g2_o21ai_1
X_4803_ _1652_ _1649_ _1657_ _1659_ VPWR VGND sg13g2_a21o_1
X_5783_ _2461_ _2463_ _2465_ _2467_ VPWR VGND sg13g2_nor3_1
X_4734_ _1601_ net488 net1496 VPWR VGND sg13g2_nand2_1
X_4665_ _1540_ _1541_ _1543_ VPWR VGND sg13g2_nor2_1
X_6404_ net556 VGND VPWR net908 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[1\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
X_3616_ _0669_ net409 _0655_ VPWR VGND sg13g2_xnor2_1
X_4596_ VGND VPWR _1480_ _1482_ _1485_ _1484_ sg13g2_a21oi_1
X_3547_ VPWR _0617_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[10\].z_sign
+ VGND sg13g2_inv_1
X_6335_ net374 _2899_ net899 _0503_ VPWR VGND sg13g2_nor3_1
X_6266_ net444 _2867_ _2868_ VPWR VGND sg13g2_and2_1
X_3478_ VPWR _0548_ net892 VGND sg13g2_inv_1
X_5217_ _1994_ net1101 _1992_ VPWR VGND sg13g2_xnor2_1
X_6197_ VGND VPWR _2808_ _2813_ _2815_ _2811_ sg13g2_a21oi_1
X_5148_ net380 VPWR _1936_ VGND _0567_ _1924_ sg13g2_o21ai_1
X_6898__549 VPWR VGND net733 sg13g2_tiehi
X_5079_ net448 net7 _0253_ VPWR VGND sg13g2_and2_1
XFILLER_13_704 VPWR VGND sg13g2_fill_1
XFILLER_5_947 VPWR VGND sg13g2_decap_8
XFILLER_47_100 VPWR VGND sg13g2_fill_2
XFILLER_0_696 VPWR VGND sg13g2_decap_8
XFILLER_48_667 VPWR VGND sg13g2_fill_2
X_6671__51 VPWR VGND net51 sg13g2_tiehi
XFILLER_28_380 VPWR VGND sg13g2_fill_2
X_6875__335 VPWR VGND net335 sg13g2_tiehi
XFILLER_11_280 VPWR VGND sg13g2_fill_1
Xhold207 _0108_ VPWR VGND net964 sg13g2_dlygate4sd3_1
X_4450_ _1362_ VPWR _1364_ VGND _1357_ _1358_ sg13g2_o21ai_1
X_4381_ _1305_ net922 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[7\]
+ VPWR VGND sg13g2_xnor2_1
Xhold229 _1378_ VPWR VGND net986 sg13g2_dlygate4sd3_1
Xhold218 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[11\] VPWR VGND net975
+ sg13g2_dlygate4sd3_1
X_6120_ _2746_ _2747_ _2748_ VPWR VGND sg13g2_nor2b_1
X_6051_ VGND VPWR _2683_ net1210 _0419_ _2688_ sg13g2_a21oi_1
X_5002_ net469 VPWR _1824_ VGND _1822_ _1823_ sg13g2_o21ai_1
X_6708__533 VPWR VGND net717 sg13g2_tiehi
XFILLER_15_0 VPWR VGND sg13g2_fill_1
XFILLER_26_339 VPWR VGND sg13g2_fill_2
X_5904_ _2562_ VPWR _2569_ VGND net512 _0576_ sg13g2_o21ai_1
X_6884_ net317 VGND VPWR _0493_ u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[4\]
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
X_5835_ net425 _2509_ _2510_ _0381_ VPWR VGND sg13g2_nor3_1
X_5766_ _2451_ _2452_ _2453_ VPWR VGND sg13g2_nor2_1
X_4717_ _1586_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[4\] _1585_
+ VPWR VGND sg13g2_nand2b_1
X_5697_ _2396_ net1519 _2395_ VPWR VGND sg13g2_nand2_1
X_6715__526 VPWR VGND net710 sg13g2_tiehi
X_4648_ _1528_ _1518_ _1524_ VPWR VGND sg13g2_nand2_1
Xhold730 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[8\] VPWR VGND net1487
+ sg13g2_dlygate4sd3_1
XFILLER_30_59 VPWR VGND sg13g2_fill_2
Xhold752 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[1\] VPWR
+ VGND net1509 sg13g2_dlygate4sd3_1
XFILLER_2_928 VPWR VGND sg13g2_decap_8
Xhold741 _2716_ VPWR VGND net1498 sg13g2_dlygate4sd3_1
Xhold763 _2406_ VPWR VGND net1520 sg13g2_dlygate4sd3_1
X_4579_ net1214 net540 _1471_ VPWR VGND sg13g2_xor2_1
Xhold796 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[5\] VPWR VGND net1553
+ sg13g2_dlygate4sd3_1
Xhold785 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[0\] VPWR
+ VGND net1542 sg13g2_dlygate4sd3_1
Xhold774 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[9\] VPWR
+ VGND net1531 sg13g2_dlygate4sd3_1
X_6318_ net465 net806 _0489_ VPWR VGND sg13g2_and2_1
X_6249_ _2855_ _2853_ _2850_ VPWR VGND sg13g2_nand2b_1
XFILLER_39_35 VPWR VGND sg13g2_fill_1
X_6722__519 VPWR VGND net703 sg13g2_tiehi
XFILLER_44_114 VPWR VGND sg13g2_fill_2
XFILLER_26_862 VPWR VGND sg13g2_fill_1
XFILLER_38_1001 VPWR VGND sg13g2_fill_2
XFILLER_5_744 VPWR VGND sg13g2_decap_8
XFILLER_4_265 VPWR VGND sg13g2_fill_2
XFILLER_20_81 VPWR VGND sg13g2_fill_1
XFILLER_49_943 VPWR VGND sg13g2_fill_2
XFILLER_1_994 VPWR VGND sg13g2_decap_8
Xhold90 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[9\] VPWR VGND net847
+ sg13g2_dlygate4sd3_1
XFILLER_35_114 VPWR VGND sg13g2_fill_2
X_3950_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[17\] u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[12\]
+ _0951_ VPWR VGND sg13g2_xor2_1
X_3881_ VGND VPWR _0537_ _0902_ _0032_ _0905_ sg13g2_a21oi_1
XFILLER_31_353 VPWR VGND sg13g2_fill_1
X_5620_ _2330_ _0598_ _2329_ VPWR VGND sg13g2_xnor2_1
X_5551_ _2268_ net934 _0338_ VPWR VGND sg13g2_nor2_1
X_4502_ VGND VPWR _1400_ _1407_ _0150_ _1408_ sg13g2_a21oi_1
X_5482_ _2213_ _2215_ _2212_ _2216_ VPWR VGND sg13g2_nand3_1
X_4433_ VGND VPWR _1350_ net387 net996 sg13g2_or2_1
Xfanout506 net939 net506 VPWR VGND sg13g2_buf_8
X_4364_ VPWR VGND _1290_ _1291_ _1280_ net411 _1292_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[7\]
+ sg13g2_a221oi_1
X_6103_ net454 VPWR _2734_ VGND _2731_ _2733_ sg13g2_o21ai_1
X_4295_ _1236_ _1232_ _1237_ VPWR VGND sg13g2_nor2b_1
Xfanout517 net518 net517 VPWR VGND sg13g2_buf_8
Xfanout528 net530 net528 VPWR VGND sg13g2_buf_8
Xfanout539 net540 net539 VPWR VGND sg13g2_buf_8
XFILLER_6_1021 VPWR VGND sg13g2_decap_8
X_6034_ _2674_ net452 _2673_ VPWR VGND sg13g2_nand2_1
XFILLER_39_431 VPWR VGND sg13g2_fill_1
XFILLER_26_125 VPWR VGND sg13g2_fill_1
XFILLER_27_659 VPWR VGND sg13g2_fill_2
X_6867_ net351 VGND VPWR _0476_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[11\]
+ clknet_leaf_7_clk sg13g2_dfrbpq_2
X_5818_ VGND VPWR _2488_ _2492_ _2495_ _2491_ sg13g2_a21oi_1
X_6798_ net627 VGND VPWR _0407_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[5\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_41_14 VPWR VGND sg13g2_fill_1
X_5749_ _2439_ net517 net1338 VPWR VGND sg13g2_nand2b_1
XFILLER_2_725 VPWR VGND sg13g2_decap_8
Xhold560 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[1\] VPWR
+ VGND net1317 sg13g2_dlygate4sd3_1
Xhold571 _0385_ VPWR VGND net1328 sg13g2_dlygate4sd3_1
Xhold582 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[3\] VPWR VGND net1339
+ sg13g2_dlygate4sd3_1
Xhold593 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[3\] VPWR VGND net1350
+ sg13g2_dlygate4sd3_1
XFILLER_1_279 VPWR VGND sg13g2_fill_2
XFILLER_32_117 VPWR VGND sg13g2_fill_2
XFILLER_12_1026 VPWR VGND sg13g2_fill_2
XFILLER_1_791 VPWR VGND sg13g2_decap_8
X_4080_ net445 _1061_ _0074_ VPWR VGND sg13g2_and2_1
X_6705__536 VPWR VGND net720 sg13g2_tiehi
X_4982_ _1798_ _1801_ _1807_ VPWR VGND sg13g2_nor2_1
X_3933_ _0935_ _0934_ net948 VPWR VGND sg13g2_nand2b_1
X_6721_ net704 VGND VPWR net1090 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[4\]
+ clknet_leaf_32_clk sg13g2_dfrbpq_1
X_3864_ VGND VPWR net842 _0890_ _0028_ _0892_ sg13g2_a21oi_1
XFILLER_31_161 VPWR VGND sg13g2_fill_1
X_6652_ net70 VGND VPWR _0261_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp\[0\]
+ clknet_leaf_16_clk sg13g2_dfrbpq_1
X_5603_ _2314_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[7\]
+ _2315_ VPWR VGND sg13g2_xor2_1
X_6583_ net139 VGND VPWR net1460 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[8\]
+ clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3795_ _0837_ _0838_ _0836_ _0842_ VPWR VGND _0841_ sg13g2_nand4_1
X_6712__529 VPWR VGND net713 sg13g2_tiehi
X_5534_ _2255_ net1507 _2257_ VPWR VGND sg13g2_and2_1
X_5465_ _2201_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[12\] _2200_
+ VPWR VGND sg13g2_xnor2_1
X_4416_ net543 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[12\] _1328_
+ _1335_ VPWR VGND sg13g2_nor3_1
X_5396_ net1386 _2132_ _2142_ VPWR VGND sg13g2_nor2_1
X_4347_ VGND VPWR _1273_ _1275_ _1278_ _1277_ sg13g2_a21oi_1
X_4278_ net497 VPWR _1222_ VGND _1217_ _1221_ sg13g2_o21ai_1
X_6017_ VGND VPWR _2652_ _2657_ _0415_ _2658_ sg13g2_a21oi_1
XFILLER_15_629 VPWR VGND sg13g2_fill_1
X_6919_ net260 VGND VPWR net960 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[13\]
+ clknet_leaf_17_clk sg13g2_dfrbpq_1
XFILLER_11_824 VPWR VGND sg13g2_fill_2
XFILLER_7_806 VPWR VGND sg13g2_decap_8
Xhold390 _2559_ VPWR VGND net1147 sg13g2_dlygate4sd3_1
XFILLER_45_220 VPWR VGND sg13g2_fill_1
XFILLER_19_968 VPWR VGND sg13g2_decap_8
XFILLER_18_456 VPWR VGND sg13g2_fill_2
XFILLER_42_993 VPWR VGND sg13g2_fill_1
XFILLER_13_161 VPWR VGND sg13g2_fill_1
XFILLER_13_194 VPWR VGND sg13g2_fill_2
X_6403__374 VPWR VGND net558 sg13g2_tiehi
X_3580_ _0633_ net860 _0001_ VPWR VGND sg13g2_nor2_1
X_5250_ _2022_ net1227 net379 VPWR VGND sg13g2_nand2_1
X_4201_ VGND VPWR _1157_ _1156_ _1151_ sg13g2_or2_1
X_5181_ net439 net913 _0275_ VPWR VGND sg13g2_nor2_1
X_4132_ VGND VPWR _1099_ _1098_ _1096_ sg13g2_or2_1
X_4063_ _0987_ _1050_ net803 _1052_ VPWR VGND sg13g2_nand3_1
XFILLER_37_743 VPWR VGND sg13g2_fill_1
X_4965_ _1792_ _1793_ _0228_ VPWR VGND sg13g2_nor2b_1
X_3916_ net463 net820 _0046_ VPWR VGND sg13g2_and2_1
X_6704_ net721 VGND VPWR _0313_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[5\]\[0\]
+ clknet_leaf_52_clk sg13g2_dfrbpq_1
X_4896_ net485 VPWR _1736_ VGND _1732_ _1734_ sg13g2_o21ai_1
X_6519__203 VPWR VGND net203 sg13g2_tiehi
X_6635_ net87 VGND VPWR net1221 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[8\]
+ clknet_leaf_24_clk sg13g2_dfrbpq_1
X_3847_ net419 net937 _0880_ _0023_ VPWR VGND sg13g2_nor3_1
X_3778_ VGND VPWR _0821_ _0823_ _0826_ _0825_ sg13g2_a21oi_1
X_6566_ net156 VGND VPWR net1213 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[4\]
+ clknet_leaf_29_clk sg13g2_dfrbpq_2
X_5517_ _2239_ _2241_ _2243_ VPWR VGND sg13g2_and2_1
X_6497_ net225 VGND VPWR net1301 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[4\]
+ clknet_leaf_32_clk sg13g2_dfrbpq_2
X_5448_ _2181_ VPWR _2186_ VGND _2178_ _2182_ sg13g2_o21ai_1
X_5379_ _2128_ _0560_ _2126_ VPWR VGND sg13g2_xnor2_1
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_47_68 VPWR VGND sg13g2_decap_8
XFILLER_15_404 VPWR VGND sg13g2_fill_1
XFILLER_16_949 VPWR VGND sg13g2_decap_8
XFILLER_24_960 VPWR VGND sg13g2_decap_8
XFILLER_23_481 VPWR VGND sg13g2_fill_1
XFILLER_11_665 VPWR VGND sg13g2_fill_2
XFILLER_7_647 VPWR VGND sg13g2_fill_1
XFILLER_3_864 VPWR VGND sg13g2_decap_8
X_6741__500 VPWR VGND net684 sg13g2_tiehi
XFILLER_18_220 VPWR VGND sg13g2_fill_1
X_6702__539 VPWR VGND net723 sg13g2_tiehi
XFILLER_18_1010 VPWR VGND sg13g2_decap_8
X_4750_ net489 VPWR _1614_ VGND _1612_ _1613_ sg13g2_o21ai_1
X_3701_ _0685_ _0636_ _0754_ VPWR VGND sg13g2_xor2_1
X_4681_ net485 VPWR _1556_ VGND _1553_ _1555_ sg13g2_o21ai_1
X_6420_ net340 VGND VPWR _0029_ u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[9\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
X_3632_ net547 u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[10\] u_angle_cordic_12b_pmod.angle_cordic_12b.COSout\[10\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[10\] net535 net545 _0685_
+ VPWR VGND sg13g2_mux4_1
X_6351_ net956 _2908_ _2911_ VPWR VGND sg13g2_nor2_1
X_3563_ net828 net445 _0528_ VPWR VGND sg13g2_and2_1
X_5302_ VGND VPWR _2058_ _2060_ _0296_ _2062_ sg13g2_a21oi_1
X_6885__315 VPWR VGND net315 sg13g2_tiehi
XFILLER_45_0 VPWR VGND sg13g2_fill_2
XFILLER_5_190 VPWR VGND sg13g2_fill_2
X_6282_ _2879_ _2868_ _0461_ VPWR VGND sg13g2_nor2b_1
X_3494_ VPWR _0564_ net529 VGND sg13g2_inv_1
X_5233_ _2008_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[12\] _1997_
+ VPWR VGND sg13g2_nand2_1
X_5164_ _1935_ VPWR _1949_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[8\]
+ net1289 sg13g2_o21ai_1
XFILLER_25_1003 VPWR VGND sg13g2_decap_8
X_4115_ _1080_ _1078_ _1083_ _1085_ VPWR VGND sg13g2_a21o_1
X_5095_ net480 VPWR _1889_ VGND _1883_ _1888_ sg13g2_o21ai_1
X_4046_ _1038_ net1012 net548 VPWR VGND sg13g2_nand2b_1
X_5997_ _2639_ _2642_ _2643_ VPWR VGND sg13g2_and2_1
X_4948_ _1779_ net1464 _1778_ VPWR VGND sg13g2_nand2_1
X_4879_ VGND VPWR _1718_ _1721_ _1719_ _1715_ sg13g2_a21oi_2
X_6618_ net104 VGND VPWR net1466 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[3\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_21_996 VPWR VGND sg13g2_decap_8
X_6549_ net173 VGND VPWR net1263 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[12\]
+ clknet_leaf_36_clk sg13g2_dfrbpq_2
XFILLER_0_801 VPWR VGND sg13g2_decap_8
XFILLER_0_878 VPWR VGND sg13g2_decap_8
XFILLER_15_223 VPWR VGND sg13g2_fill_2
XFILLER_8_923 VPWR VGND sg13g2_decap_8
XFILLER_12_963 VPWR VGND sg13g2_decap_8
XFILLER_48_1014 VPWR VGND sg13g2_decap_8
X_6509__213 VPWR VGND net213 sg13g2_tiehi
XFILLER_38_348 VPWR VGND sg13g2_fill_1
X_5920_ VGND VPWR _0579_ _2575_ _2583_ net512 sg13g2_a21oi_1
X_5851_ VGND VPWR _2519_ net1347 _0383_ _2524_ sg13g2_a21oi_1
X_4802_ _1652_ _1657_ _1649_ _1658_ VPWR VGND sg13g2_nand3_1
X_5782_ _2465_ VPWR _2466_ VGND _2461_ _2463_ sg13g2_o21ai_1
X_4733_ _1593_ _1597_ _1598_ _1600_ VPWR VGND sg13g2_nor3_1
X_6516__206 VPWR VGND net206 sg13g2_tiehi
X_6403_ net558 VGND VPWR net884 u_angle_cordic_12b_pmod.u_vga_top.v_pos\[0\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
X_4664_ _1540_ _1541_ _1542_ VPWR VGND sg13g2_and2_1
X_3615_ VPWR _0668_ _0667_ VGND sg13g2_inv_1
X_4595_ net1185 net540 _1484_ VPWR VGND sg13g2_xor2_1
X_3546_ VPWR _0616_ net1556 VGND sg13g2_inv_1
X_6334_ net898 _2898_ _2900_ VPWR VGND sg13g2_nor2_1
X_6265_ net1041 VPWR _2867_ VGND net967 net555 sg13g2_o21ai_1
X_5216_ net1101 _1992_ _1993_ VPWR VGND sg13g2_nor2_1
X_3477_ VPWR _0547_ net1107 VGND sg13g2_inv_1
X_6196_ VGND VPWR _2807_ net1344 _0438_ _2814_ sg13g2_a21oi_1
X_5147_ VPWR _1935_ net380 VGND sg13g2_inv_1
XFILLER_28_37 VPWR VGND sg13g2_fill_1
X_5078_ net448 net6 _0252_ VPWR VGND sg13g2_and2_1
X_4029_ _1018_ VPWR _1024_ VGND _1016_ _1017_ sg13g2_o21ai_1
XFILLER_37_370 VPWR VGND sg13g2_fill_1
XFILLER_8_219 VPWR VGND sg13g2_fill_2
X_6731__510 VPWR VGND net694 sg13g2_tiehi
XFILLER_5_926 VPWR VGND sg13g2_decap_8
XFILLER_0_642 VPWR VGND sg13g2_fill_1
XFILLER_47_112 VPWR VGND sg13g2_fill_1
XFILLER_0_675 VPWR VGND sg13g2_decap_8
XFILLER_16_576 VPWR VGND sg13g2_decap_4
Xhold208 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[1\] VPWR VGND net965
+ sg13g2_dlygate4sd3_1
Xhold219 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[0\] VPWR VGND net976
+ sg13g2_dlygate4sd3_1
X_4380_ net922 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[7\] _1304_
+ VPWR VGND sg13g2_nor2b_1
X_6050_ net452 VPWR _2688_ VGND _2683_ _2687_ sg13g2_o21ai_1
XFILLER_22_2 VPWR VGND sg13g2_fill_1
X_5001_ _1823_ net1196 net399 VPWR VGND sg13g2_xnor2_1
XFILLER_22_1028 VPWR VGND sg13g2_fill_1
X_6883_ net319 VGND VPWR _0492_ u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[3\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_1
X_5903_ _2565_ _2561_ _2564_ _2568_ VPWR VGND sg13g2_a21o_1
X_5834_ _2508_ _2503_ _2510_ VPWR VGND sg13g2_nor2b_1
X_5765_ VGND VPWR _2446_ _2447_ _2452_ _2448_ sg13g2_a21oi_1
X_4716_ _1585_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[10\]
+ _1584_ VPWR VGND sg13g2_xnor2_1
X_5696_ _2395_ net1467 _2394_ VPWR VGND sg13g2_xnor2_1
X_4647_ net432 _1526_ _1527_ _0176_ VPWR VGND sg13g2_nor3_1
XFILLER_2_907 VPWR VGND sg13g2_decap_8
Xhold720 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[8\] VPWR VGND net1477
+ sg13g2_dlygate4sd3_1
Xhold731 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[2\] VPWR VGND net1488
+ sg13g2_dlygate4sd3_1
X_6317_ VGND VPWR _0605_ net815 _0488_ _2897_ sg13g2_a21oi_1
Xhold753 _2572_ VPWR VGND net1510 sg13g2_dlygate4sd3_1
Xhold764 _0359_ VPWR VGND net1521 sg13g2_dlygate4sd3_1
Xhold742 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[6\]\[4\] VPWR VGND net1499
+ sg13g2_dlygate4sd3_1
X_4578_ _1470_ _0608_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[8\]\[6\]
+ VPWR VGND sg13g2_nand2_1
Xhold797 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[5\] VPWR
+ VGND net1554 sg13g2_dlygate4sd3_1
X_3529_ VPWR _0599_ net1482 VGND sg13g2_inv_1
Xhold786 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[10\]\[4\] VPWR VGND net1543
+ sg13g2_dlygate4sd3_1
Xhold775 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[9\] VPWR VGND net1532
+ sg13g2_dlygate4sd3_1
X_6248_ VGND VPWR _2852_ _2853_ _0450_ _2854_ sg13g2_a21oi_1
X_6179_ VGND VPWR _2793_ _2798_ _0436_ _2799_ sg13g2_a21oi_1
XFILLER_13_513 VPWR VGND sg13g2_fill_2
XFILLER_5_723 VPWR VGND sg13g2_decap_8
XFILLER_1_973 VPWR VGND sg13g2_decap_8
X_6629__93 VPWR VGND net93 sg13g2_tiehi
Xhold80 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[10\] VPWR VGND net837
+ sg13g2_dlygate4sd3_1
Xhold91 _0510_ VPWR VGND net848 sg13g2_dlygate4sd3_1
X_6506__216 VPWR VGND net216 sg13g2_tiehi
X_3880_ net443 VPWR _0905_ VGND _0537_ _0902_ sg13g2_o21ai_1
XFILLER_31_332 VPWR VGND sg13g2_fill_1
X_5550_ net474 VPWR _2269_ VGND net933 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[0\]
+ sg13g2_o21ai_1
X_4501_ net489 VPWR _1408_ VGND _1400_ _1407_ sg13g2_o21ai_1
X_5481_ VPWR _2215_ _2214_ VGND sg13g2_inv_1
X_4432_ _1349_ net996 net386 VPWR VGND sg13g2_nand2_1
X_6513__209 VPWR VGND net209 sg13g2_tiehi
X_4363_ _1291_ _1283_ _1281_ VPWR VGND sg13g2_nand2b_1
X_6413__354 VPWR VGND net354 sg13g2_tiehi
Xfanout507 net511 net507 VPWR VGND sg13g2_buf_8
X_6102_ _2732_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[12\] _2733_
+ VPWR VGND sg13g2_xor2_1
X_4294_ _1236_ net1462 net381 VPWR VGND sg13g2_xnor2_1
Xfanout518 net519 net518 VPWR VGND sg13g2_buf_8
Xfanout529 net530 net529 VPWR VGND sg13g2_buf_1
XFILLER_6_1000 VPWR VGND sg13g2_decap_8
X_6033_ VGND VPWR _2673_ _2672_ _2667_ sg13g2_or2_1
XFILLER_27_627 VPWR VGND sg13g2_fill_1
X_6721__520 VPWR VGND net704 sg13g2_tiehi
XFILLER_23_800 VPWR VGND sg13g2_fill_1
XFILLER_41_129 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_61_clk clknet_4_2_0_clk clknet_leaf_61_clk VPWR VGND sg13g2_buf_8
X_6866_ net353 VGND VPWR _0475_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[10\]
+ clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_34_192 VPWR VGND sg13g2_fill_1
X_5817_ VGND VPWR _2488_ _2493_ _0379_ _2494_ sg13g2_a21oi_1
X_6797_ net628 VGND VPWR _0406_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[4\]
+ clknet_leaf_10_clk sg13g2_dfrbpq_1
X_5748_ net517 net1338 _2438_ VPWR VGND sg13g2_nor2b_1
X_5679_ net412 _2373_ _2380_ VPWR VGND sg13g2_and2_1
XFILLER_2_704 VPWR VGND sg13g2_decap_8
Xhold550 _2516_ VPWR VGND net1307 sg13g2_dlygate4sd3_1
Xhold561 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[7\] VPWR VGND net1318
+ sg13g2_dlygate4sd3_1
Xhold572 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[4\] VPWR VGND net1329
+ sg13g2_dlygate4sd3_1
Xhold594 _1510_ VPWR VGND net1351 sg13g2_dlygate4sd3_1
Xhold583 _0417_ VPWR VGND net1340 sg13g2_dlygate4sd3_1
XFILLER_46_925 VPWR VGND sg13g2_fill_2
X_6626__96 VPWR VGND net96 sg13g2_tiehi
X_6837__404 VPWR VGND net588 sg13g2_tiehi
Xclkbuf_leaf_52_clk clknet_4_10_0_clk clknet_leaf_52_clk VPWR VGND sg13g2_buf_8
XFILLER_13_376 VPWR VGND sg13g2_fill_1
XFILLER_14_899 VPWR VGND sg13g2_decap_8
XFILLER_12_1005 VPWR VGND sg13g2_decap_8
XFILLER_1_770 VPWR VGND sg13g2_decap_8
XFILLER_49_752 VPWR VGND sg13g2_fill_1
X_4981_ VGND VPWR _1804_ _1805_ _0231_ _1806_ sg13g2_a21oi_1
X_3932_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[2\] _0933_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[3\]
+ _0934_ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_43_clk clknet_4_14_0_clk clknet_leaf_43_clk VPWR VGND sg13g2_buf_8
X_6720_ net705 VGND VPWR _0329_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[3\]
+ clknet_leaf_30_clk sg13g2_dfrbpq_2
X_6651_ net71 VGND VPWR _0260_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[12\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_1
X_3863_ _0885_ VPWR _0892_ VGND net842 _0890_ sg13g2_o21ai_1
X_6582_ net140 VGND VPWR _0191_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[7\]
+ clknet_leaf_34_clk sg13g2_dfrbpq_2
X_5602_ net516 _2313_ _2314_ VPWR VGND sg13g2_nor2_1
X_3794_ net863 net813 _0839_ _0840_ _0841_ VPWR VGND sg13g2_nor4_1
X_5533_ net418 VPWR _2256_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[6\]
+ net1156 sg13g2_o21ai_1
X_5464_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[11\] net418 _2194_
+ _2200_ VPWR VGND sg13g2_a21o_1
X_5395_ VGND VPWR _2137_ _2139_ _2141_ _2136_ sg13g2_a21oi_1
X_4415_ VGND VPWR _1326_ _1331_ _1334_ _1330_ sg13g2_a21oi_1
X_4346_ net1120 net541 _1277_ VPWR VGND sg13g2_xor2_1
X_4277_ _1221_ net1404 _1219_ VPWR VGND sg13g2_xnor2_1
X_6016_ net452 VPWR _2658_ VGND _2652_ _2657_ sg13g2_o21ai_1
XFILLER_36_48 VPWR VGND sg13g2_fill_1
XFILLER_14_118 VPWR VGND sg13g2_fill_1
X_6623__99 VPWR VGND net99 sg13g2_tiehi
Xclkbuf_leaf_34_clk clknet_4_13_0_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
X_6918_ net262 VGND VPWR _0513_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[12\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
X_6849_ net576 VGND VPWR _0458_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[6\]
+ clknet_leaf_63_clk sg13g2_dfrbpq_2
XFILLER_2_545 VPWR VGND sg13g2_fill_2
Xhold380 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[8\] VPWR VGND net1137
+ sg13g2_dlygate4sd3_1
Xhold391 _0390_ VPWR VGND net1148 sg13g2_dlygate4sd3_1
XFILLER_2_578 VPWR VGND sg13g2_fill_1
XFILLER_46_722 VPWR VGND sg13g2_fill_2
XFILLER_19_947 VPWR VGND sg13g2_decap_8
X_6503__219 VPWR VGND net219 sg13g2_tiehi
Xclkbuf_leaf_25_clk clknet_4_13_0_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
XFILLER_10_880 VPWR VGND sg13g2_decap_8
X_6711__530 VPWR VGND net714 sg13g2_tiehi
XFILLER_6_895 VPWR VGND sg13g2_decap_8
X_4200_ _1156_ net991 _1154_ VPWR VGND sg13g2_xnor2_1
X_5180_ _1962_ net912 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[5\]
+ VPWR VGND sg13g2_xnor2_1
X_4131_ net1175 net533 _1098_ VPWR VGND sg13g2_xor2_1
X_4062_ VGND VPWR _0992_ _1050_ _1051_ _0082_ sg13g2_a21oi_1
XFILLER_37_700 VPWR VGND sg13g2_fill_2
XFILLER_3_1025 VPWR VGND sg13g2_decap_4
X_4964_ net469 _1791_ _1793_ VPWR VGND sg13g2_and2_1
Xclkbuf_leaf_16_clk clknet_4_4_0_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
X_6703_ net722 VGND VPWR net1234 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[12\]
+ clknet_leaf_56_clk sg13g2_dfrbpq_2
X_3915_ net463 net790 _0045_ VPWR VGND sg13g2_and2_1
X_4895_ _1735_ _1732_ _1734_ VPWR VGND sg13g2_nand2_1
X_6634_ net88 VGND VPWR net1431 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[7\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_1
X_3846_ net936 _0878_ _0880_ VPWR VGND sg13g2_and2_1
X_3777_ net978 net920 net1024 _0824_ _0825_ VPWR VGND sg13g2_nor4_1
X_6565_ net157 VGND VPWR net1353 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[3\]
+ clknet_leaf_26_clk sg13g2_dfrbpq_1
X_6496_ net226 VGND VPWR _0105_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[3\]
+ clknet_leaf_46_clk sg13g2_dfrbpq_2
X_5516_ VGND VPWR _2238_ _2240_ _0330_ _2242_ sg13g2_a21oi_1
X_5447_ net429 _2184_ _2185_ _0318_ VPWR VGND sg13g2_nor3_1
X_6391__541 VPWR VGND net725 sg13g2_tiehi
X_5378_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[8\] _2126_ _2127_
+ VPWR VGND sg13g2_and2_1
X_6827__414 VPWR VGND net598 sg13g2_tiehi
X_4329_ VGND VPWR net770 _1261_ _1263_ _1260_ sg13g2_a21oi_1
XFILLER_16_928 VPWR VGND sg13g2_decap_8
X_6834__407 VPWR VGND net591 sg13g2_tiehi
XFILLER_11_655 VPWR VGND sg13g2_fill_2
XFILLER_3_843 VPWR VGND sg13g2_decap_8
XFILLER_21_408 VPWR VGND sg13g2_fill_1
XFILLER_15_983 VPWR VGND sg13g2_decap_8
X_3700_ _0753_ _0636_ _0685_ VPWR VGND sg13g2_nand2_1
X_4680_ _1555_ net1177 net394 VPWR VGND sg13g2_xnor2_1
X_3631_ VPWR _0684_ _0683_ VGND sg13g2_inv_1
X_3562_ _0531_ net422 _0527_ VPWR VGND sg13g2_nor2_1
X_6350_ net956 _2908_ _2910_ VPWR VGND sg13g2_and2_1
X_5301_ _2062_ net497 _2061_ VPWR VGND sg13g2_nand2_1
X_6281_ net421 _2873_ _2880_ _0460_ VPWR VGND sg13g2_nor3_1
X_3493_ VPWR _0563_ net1392 VGND sg13g2_inv_1
X_5232_ VGND VPWR _2006_ _2007_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[12\]
+ net526 sg13g2_a21oi_2
Xclkbuf_leaf_5_clk clknet_4_1_0_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_5163_ _1941_ _1944_ _1940_ _1948_ VPWR VGND sg13g2_nand3_1
X_4114_ _1080_ _1083_ _1078_ _1084_ VPWR VGND sg13g2_nand3_1
X_5094_ _1888_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[1\] _1886_
+ VPWR VGND sg13g2_xnor2_1
XFILLER_37_552 VPWR VGND sg13g2_fill_1
X_4045_ _1037_ _0939_ _1034_ VPWR VGND sg13g2_nand2_1
XFILLER_24_202 VPWR VGND sg13g2_fill_1
XFILLER_13_909 VPWR VGND sg13g2_decap_8
XFILLER_25_736 VPWR VGND sg13g2_fill_1
XFILLER_24_257 VPWR VGND sg13g2_fill_1
X_5996_ _0410_ net460 _2641_ _2642_ VPWR VGND sg13g2_and3_1
X_4947_ _1777_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[12\] _1778_
+ VPWR VGND sg13g2_xor2_1
X_4878_ VGND VPWR _1715_ _1719_ _0214_ _1720_ sg13g2_a21oi_1
XFILLER_21_975 VPWR VGND sg13g2_decap_8
X_6617_ net105 VGND VPWR _0226_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[2\]
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
X_3829_ net553 net869 _0868_ VPWR VGND sg13g2_nor2_1
X_6548_ net174 VGND VPWR net1170 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[11\]
+ clknet_leaf_37_clk sg13g2_dfrbpq_2
X_6479_ net243 VGND VPWR net1061 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[5\]
+ clknet_leaf_42_clk sg13g2_dfrbpq_1
XFILLER_0_857 VPWR VGND sg13g2_decap_8
X_6701__540 VPWR VGND net724 sg13g2_tiehi
XFILLER_43_588 VPWR VGND sg13g2_fill_2
XFILLER_8_902 VPWR VGND sg13g2_decap_8
XFILLER_12_942 VPWR VGND sg13g2_decap_8
XFILLER_8_979 VPWR VGND sg13g2_decap_8
XFILLER_7_467 VPWR VGND sg13g2_fill_1
XFILLER_7_434 VPWR VGND sg13g2_fill_1
XFILLER_3_640 VPWR VGND sg13g2_fill_2
XFILLER_47_850 VPWR VGND sg13g2_fill_1
X_5850_ net458 VPWR _2524_ VGND _2519_ _2523_ sg13g2_o21ai_1
X_6817__424 VPWR VGND net608 sg13g2_tiehi
X_5781_ _2465_ net520 net1127 VPWR VGND sg13g2_xnor2_1
X_4801_ _1657_ net1383 _1655_ VPWR VGND sg13g2_xnor2_1
X_4732_ _1597_ VPWR _1599_ VGND _1593_ _1598_ sg13g2_o21ai_1
XFILLER_14_290 VPWR VGND sg13g2_fill_2
X_4663_ _1541_ net1017 net393 VPWR VGND sg13g2_xnor2_1
X_3614_ _0667_ net409 _0655_ VPWR VGND sg13g2_nand2_1
X_6402_ net559 VGND VPWR _0011_ pwm_data clknet_leaf_13_clk sg13g2_dfrbpq_1
X_4594_ VGND VPWR _1479_ net1087 _0167_ _1483_ sg13g2_a21oi_1
X_3545_ VPWR _0615_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[2\]
+ VGND sg13g2_inv_1
X_6333_ net898 _2898_ _2899_ VPWR VGND sg13g2_and2_1
X_6264_ _2864_ _2865_ _2866_ VPWR VGND sg13g2_nor2b_1
X_3476_ VPWR _0546_ net459 VGND sg13g2_inv_1
X_5215_ _1992_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[10\] _1991_
+ VPWR VGND sg13g2_xnor2_1
X_6824__417 VPWR VGND net601 sg13g2_tiehi
X_6195_ net454 VPWR _2814_ VGND _2807_ _2812_ sg13g2_o21ai_1
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk VPWR VGND sg13g2_buf_8
X_5146_ VGND VPWR _1932_ _1934_ _1933_ _1924_ sg13g2_a21oi_2
X_5077_ net448 net5 _0251_ VPWR VGND sg13g2_and2_1
X_6680__42 VPWR VGND net42 sg13g2_tiehi
X_4028_ _1023_ net952 net549 VPWR VGND sg13g2_xnor2_1
X_6423__334 VPWR VGND net334 sg13g2_tiehi
X_5979_ net467 net783 _0405_ VPWR VGND sg13g2_and2_1
XFILLER_5_905 VPWR VGND sg13g2_decap_8
XFILLER_0_654 VPWR VGND sg13g2_decap_8
XFILLER_47_102 VPWR VGND sg13g2_fill_1
XFILLER_48_669 VPWR VGND sg13g2_fill_1
XFILLER_48_647 VPWR VGND sg13g2_fill_1
X_6467__261 VPWR VGND net261 sg13g2_tiehi
XFILLER_16_522 VPWR VGND sg13g2_fill_1
XFILLER_18_93 VPWR VGND sg13g2_fill_2
XFILLER_15_1025 VPWR VGND sg13g2_decap_4
Xhold209 _2736_ VPWR VGND net966 sg13g2_dlygate4sd3_1
XFILLER_4_993 VPWR VGND sg13g2_decap_8
X_5000_ VGND VPWR net1052 net399 _1822_ _1821_ sg13g2_a21oi_1
XFILLER_22_1007 VPWR VGND sg13g2_decap_8
X_6446__301 VPWR VGND net301 sg13g2_tiehi
XFILLER_38_146 VPWR VGND sg13g2_fill_2
X_6522__200 VPWR VGND net200 sg13g2_tiehi
X_6882_ net321 VGND VPWR _0491_ u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[2\]
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
X_5902_ _2566_ _2567_ _0391_ VPWR VGND sg13g2_nor2b_1
X_5833_ _2503_ _2508_ _2509_ VPWR VGND sg13g2_nor2b_1
X_5764_ _2451_ net518 net1354 VPWR VGND sg13g2_xnor2_1
X_4715_ net537 _1558_ _1584_ VPWR VGND sg13g2_nor2_1
X_5695_ VGND VPWR _0599_ _2386_ _2394_ net516 sg13g2_a21oi_1
X_4646_ _1527_ _1518_ _1520_ _1525_ VPWR VGND sg13g2_and3_1
X_4577_ _1467_ _1468_ _1469_ VPWR VGND sg13g2_nor2_1
Xhold721 _0155_ VPWR VGND net1478 sg13g2_dlygate4sd3_1
Xhold710 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[10\] VPWR VGND net1467
+ sg13g2_dlygate4sd3_1
Xhold743 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[3\] VPWR VGND net1500
+ sg13g2_dlygate4sd3_1
Xhold732 _1839_ VPWR VGND net1489 sg13g2_dlygate4sd3_1
Xhold754 _0392_ VPWR VGND net1511 sg13g2_dlygate4sd3_1
X_6316_ _2896_ _2897_ _0487_ VPWR VGND sg13g2_nor2_1
Xhold776 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[5\] VPWR VGND net1533
+ sg13g2_dlygate4sd3_1
Xhold765 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[6\] VPWR VGND net1522
+ sg13g2_dlygate4sd3_1
X_3528_ _0598_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[10\]
+ VPWR VGND sg13g2_inv_2
Xhold787 _1799_ VPWR VGND net1544 sg13g2_dlygate4sd3_1
Xhold798 _0396_ VPWR VGND net1555 sg13g2_dlygate4sd3_1
X_6247_ net455 VPWR _2854_ VGND _2852_ _2853_ sg13g2_o21ai_1
X_6178_ net454 VPWR _2799_ VGND _2793_ _2798_ sg13g2_o21ai_1
X_5129_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[5\] _1918_ _1919_
+ VPWR VGND sg13g2_nor2_1
XFILLER_44_116 VPWR VGND sg13g2_fill_1
XFILLER_40_377 VPWR VGND sg13g2_fill_1
XFILLER_21_580 VPWR VGND sg13g2_fill_1
XFILLER_5_779 VPWR VGND sg13g2_decap_8
XFILLER_1_952 VPWR VGND sg13g2_decap_8
X_6807__434 VPWR VGND net618 sg13g2_tiehi
XFILLER_48_422 VPWR VGND sg13g2_fill_1
Xhold70 _0375_ VPWR VGND net827 sg13g2_dlygate4sd3_1
Xhold81 _0299_ VPWR VGND net838 sg13g2_dlygate4sd3_1
Xhold92 u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[3\] VPWR VGND net849 sg13g2_dlygate4sd3_1
XFILLER_35_116 VPWR VGND sg13g2_fill_1
XFILLER_44_661 VPWR VGND sg13g2_fill_1
X_6814__427 VPWR VGND net611 sg13g2_tiehi
X_5480_ _2202_ VPWR _2214_ VGND _0557_ _2206_ sg13g2_o21ai_1
X_4500_ _1407_ net1442 _1405_ VPWR VGND sg13g2_nand2b_1
X_4431_ _1348_ _1347_ _1343_ VPWR VGND sg13g2_nand2b_1
X_4362_ _1284_ _1287_ _1290_ VPWR VGND sg13g2_nor2_1
XFILLER_4_790 VPWR VGND sg13g2_decap_8
X_6101_ _2724_ net510 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[11\]
+ _2732_ VPWR VGND sg13g2_mux2_1
X_4293_ net381 net1567 _1235_ VPWR VGND sg13g2_nor2b_1
Xfanout508 net509 net508 VPWR VGND sg13g2_buf_8
Xfanout519 net520 net519 VPWR VGND sg13g2_buf_8
X_6032_ _2672_ net1339 _2670_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_0 VPWR VGND sg13g2_fill_2
X_6865_ net355 VGND VPWR _0474_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[9\]
+ clknet_leaf_7_clk sg13g2_dfrbpq_2
X_5816_ net457 VPWR _2494_ VGND _2488_ _2493_ sg13g2_o21ai_1
XFILLER_23_878 VPWR VGND sg13g2_fill_2
X_6796_ net629 VGND VPWR _0405_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[3\]
+ clknet_leaf_29_clk sg13g2_dfrbpq_1
X_5747_ _2434_ VPWR _2437_ VGND _2433_ _2435_ sg13g2_o21ai_1
X_5678_ VGND VPWR _2371_ _2376_ _2379_ _2375_ sg13g2_a21oi_1
X_4629_ _1506_ _1510_ _1512_ VPWR VGND sg13g2_nor2b_1
Xhold551 _0382_ VPWR VGND net1308 sg13g2_dlygate4sd3_1
Xhold540 _0418_ VPWR VGND net1297 sg13g2_dlygate4sd3_1
Xhold562 _2700_ VPWR VGND net1319 sg13g2_dlygate4sd3_1
Xhold584 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[11\] VPWR VGND net1341
+ sg13g2_dlygate4sd3_1
Xhold595 _1511_ VPWR VGND net1352 sg13g2_dlygate4sd3_1
Xhold573 _2833_ VPWR VGND net1330 sg13g2_dlygate4sd3_1
XFILLER_41_620 VPWR VGND sg13g2_fill_2
XFILLER_14_878 VPWR VGND sg13g2_decap_8
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
X_6436__311 VPWR VGND net311 sg13g2_tiehi
X_6512__210 VPWR VGND net210 sg13g2_tiehi
X_6443__304 VPWR VGND net304 sg13g2_tiehi
XFILLER_23_108 VPWR VGND sg13g2_fill_2
X_4980_ net467 VPWR _1806_ VGND _1804_ _1805_ sg13g2_o21ai_1
X_3931_ VGND VPWR _0933_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[0\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[1\] sg13g2_or2_1
XFILLER_17_694 VPWR VGND sg13g2_fill_2
X_3862_ _0890_ net1020 _0027_ VPWR VGND sg13g2_nor2_1
X_6650_ net72 VGND VPWR _0259_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg\[11\]
+ clknet_leaf_18_clk sg13g2_dfrbpq_1
X_6581_ net141 VGND VPWR _0190_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[6\]
+ clknet_leaf_34_clk sg13g2_dfrbpq_2
X_5601_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[5\] u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[6\]
+ _2295_ _2313_ VPWR VGND sg13g2_nor3_1
X_3793_ net866 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[6\] _0840_ VPWR VGND sg13g2_xor2_1
X_5532_ _2255_ _2253_ _2251_ VPWR VGND sg13g2_nand2b_1
X_5463_ _2196_ VPWR _2199_ VGND _2193_ _2197_ sg13g2_o21ai_1
X_5394_ VGND VPWR _2137_ _2139_ _0310_ _2140_ sg13g2_a21oi_1
X_4414_ net1375 _1333_ _0137_ VPWR VGND sg13g2_nor2b_1
XFILLER_28_1013 VPWR VGND sg13g2_decap_8
X_4345_ VGND VPWR _1272_ _1274_ _0125_ _1276_ sg13g2_a21oi_1
X_4276_ _1220_ net1404 _1219_ VPWR VGND sg13g2_nand2_1
X_6015_ _2657_ _0545_ _2655_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_414 VPWR VGND sg13g2_fill_2
X_6917_ net264 VGND VPWR _0512_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[11\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
X_6848_ net577 VGND VPWR _0457_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[5\]
+ clknet_leaf_63_clk sg13g2_dfrbpq_2
XFILLER_11_826 VPWR VGND sg13g2_fill_1
X_6779_ net646 VGND VPWR net1218 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[12\]
+ clknet_leaf_58_clk sg13g2_dfrbpq_2
Xhold370 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[9\] VPWR VGND net1127
+ sg13g2_dlygate4sd3_1
Xhold381 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[7\] VPWR VGND net1138
+ sg13g2_dlygate4sd3_1
Xhold392 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[8\] VPWR VGND net1149
+ sg13g2_dlygate4sd3_1
XFILLER_18_414 VPWR VGND sg13g2_fill_1
XFILLER_19_926 VPWR VGND sg13g2_decap_8
X_6804__437 VPWR VGND net621 sg13g2_tiehi
XFILLER_18_458 VPWR VGND sg13g2_fill_1
XFILLER_27_981 VPWR VGND sg13g2_decap_8
XFILLER_6_874 VPWR VGND sg13g2_decap_8
X_4130_ _1097_ _0582_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[7\]
+ VPWR VGND sg13g2_nand2_1
X_4061_ _1049_ VPWR _1050_ VGND _1045_ _1046_ sg13g2_o21ai_1
XFILLER_3_1004 VPWR VGND sg13g2_decap_8
X_4963_ VGND VPWR _1788_ _1789_ _1792_ _1790_ sg13g2_a21oi_1
X_3914_ net464 net774 _0044_ VPWR VGND sg13g2_and2_1
X_6702_ net723 VGND VPWR net1387 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[11\]
+ clknet_leaf_49_clk sg13g2_dfrbpq_2
X_4894_ net389 net1251 _1734_ VPWR VGND sg13g2_xor2_1
X_6633_ net89 VGND VPWR net1561 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[6\]
+ clknet_leaf_19_clk sg13g2_dfrbpq_1
XFILLER_32_472 VPWR VGND sg13g2_fill_1
X_3845_ net936 _0878_ _0879_ VPWR VGND sg13g2_nor2_1
X_6564_ net158 VGND VPWR _0173_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[2\]
+ clknet_leaf_36_clk sg13g2_dfrbpq_2
X_3776_ net941 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[5\] u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[7\]
+ _0824_ VPWR VGND u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[4\] sg13g2_nand4_1
X_6495_ net227 VGND VPWR net1184 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[2\]
+ clknet_leaf_45_clk sg13g2_dfrbpq_2
X_5515_ _2242_ net481 _2241_ VPWR VGND sg13g2_nand2_1
X_5446_ _2178_ _2183_ _2185_ VPWR VGND sg13g2_nor2b_1
X_6454__285 VPWR VGND net285 sg13g2_tiehi
X_5377_ _2125_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[10\]
+ _2126_ VPWR VGND sg13g2_xor2_1
X_4328_ VGND VPWR net770 _1261_ _0122_ _1262_ sg13g2_a21oi_1
XFILLER_47_15 VPWR VGND sg13g2_decap_4
X_4259_ _1205_ net1322 _1203_ VPWR VGND sg13g2_xnor2_1
XFILLER_16_907 VPWR VGND sg13g2_decap_8
XFILLER_15_439 VPWR VGND sg13g2_fill_2
X_6502__220 VPWR VGND net220 sg13g2_tiehi
XFILLER_24_995 VPWR VGND sg13g2_decap_8
XFILLER_3_822 VPWR VGND sg13g2_decap_8
X_6433__314 VPWR VGND net314 sg13g2_tiehi
XFILLER_3_899 VPWR VGND sg13g2_decap_8
XFILLER_2_376 VPWR VGND sg13g2_fill_2
XFILLER_2_387 VPWR VGND sg13g2_fill_1
X_6440__307 VPWR VGND net307 sg13g2_tiehi
XFILLER_15_962 VPWR VGND sg13g2_decap_8
X_6618__104 VPWR VGND net104 sg13g2_tiehi
X_3630_ _0655_ net405 _0682_ _0683_ VPWR VGND sg13g2_a21o_1
X_3561_ net824 net445 _0526_ VPWR VGND sg13g2_and2_1
X_5300_ VGND VPWR _2061_ _2060_ _2058_ sg13g2_or2_1
X_6280_ VPWR VGND net1041 _2864_ _2876_ net939 _2880_ net1070 sg13g2_a221oi_1
X_3492_ VPWR _0562_ net509 VGND sg13g2_inv_1
X_5231_ net526 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[12\] _1997_
+ _2006_ VPWR VGND sg13g2_nor3_1
X_5162_ _1947_ _0571_ net380 VPWR VGND sg13g2_xnor2_1
X_5093_ _1887_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[1\] _1886_
+ VPWR VGND sg13g2_nand2_1
X_4113_ net1266 net532 _1083_ VPWR VGND sg13g2_xor2_1
X_4044_ _1031_ VPWR _0064_ VGND _1035_ _1036_ sg13g2_o21ai_1
X_5995_ _2637_ _2635_ _2640_ _2642_ VPWR VGND sg13g2_a21o_1
X_4946_ _0617_ VPWR _1777_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[10\]
+ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[11\] sg13g2_o21ai_1
XFILLER_21_910 VPWR VGND sg13g2_fill_2
X_4877_ net483 VPWR _1720_ VGND _1715_ _1719_ sg13g2_o21ai_1
XFILLER_21_954 VPWR VGND sg13g2_decap_8
X_6616_ net106 VGND VPWR net1161 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[1\]
+ clknet_leaf_23_clk sg13g2_dfrbpq_1
X_3828_ net867 _0867_ _0017_ VPWR VGND sg13g2_nor2b_1
X_6547_ net175 VGND VPWR _0156_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[10\]
+ clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3759_ _0811_ VPWR _0812_ VGND _0788_ _0799_ sg13g2_o21ai_1
X_6478_ net244 VGND VPWR _0087_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[4\]
+ clknet_leaf_42_clk sg13g2_dfrbpq_1
X_5429_ net477 VPWR _2170_ VGND _2164_ _2169_ sg13g2_o21ai_1
XFILLER_0_836 VPWR VGND sg13g2_decap_8
X_6840__401 VPWR VGND net585 sg13g2_tiehi
XFILLER_15_225 VPWR VGND sg13g2_fill_1
XFILLER_12_921 VPWR VGND sg13g2_decap_8
XFILLER_12_998 VPWR VGND sg13g2_decap_8
XFILLER_8_958 VPWR VGND sg13g2_decap_8
X_6400__379 VPWR VGND net563 sg13g2_tiehi
XFILLER_3_696 VPWR VGND sg13g2_decap_8
XFILLER_48_91 VPWR VGND sg13g2_fill_1
XFILLER_0_1018 VPWR VGND sg13g2_decap_8
XFILLER_0_76 VPWR VGND sg13g2_fill_2
X_4800_ _1656_ net1383 _1655_ VPWR VGND sg13g2_nand2_1
X_5780_ _2463_ _2464_ _0372_ VPWR VGND sg13g2_nor2b_1
X_4731_ VPWR VGND net1293 _1587_ net401 _1583_ _1598_ _1588_ sg13g2_a221oi_1
X_4662_ VPWR VGND _1538_ _1539_ _1529_ net1189 _1540_ net393 sg13g2_a221oi_1
X_6401_ net561 VGND VPWR net1067 net22 clknet_leaf_0_clk sg13g2_dfrbpq_1
X_3613_ VGND VPWR _0664_ _0665_ _0666_ _0659_ sg13g2_a21oi_1
XFILLER_31_1020 VPWR VGND sg13g2_decap_8
X_4593_ _1483_ net503 _1482_ VPWR VGND sg13g2_nand2_1
X_6332_ _0958_ net374 _2898_ _0502_ VPWR VGND sg13g2_nor3_1
X_6889__294 VPWR VGND net294 sg13g2_tiehi
X_3544_ VPWR _0614_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[1\] VGND
+ sg13g2_inv_1
X_6263_ net1070 VPWR _2865_ VGND net506 _2863_ sg13g2_o21ai_1
X_3475_ VPWR _0545_ net965 VGND sg13g2_inv_1
X_5214_ VGND VPWR _0570_ _1984_ _1991_ net527 sg13g2_a21oi_1
X_6194_ VPWR _2813_ _2812_ VGND sg13g2_inv_1
X_5145_ net527 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[10\]
+ _1933_ VPWR VGND sg13g2_nor2_1
X_5076_ net448 net4 _0250_ VPWR VGND sg13g2_and2_1
X_4027_ net549 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[6\] _1022_
+ VPWR VGND sg13g2_nor2b_1
X_5978_ net467 net766 _0404_ VPWR VGND sg13g2_and2_1
X_4929_ VGND VPWR _1761_ _1762_ _0222_ _1763_ sg13g2_a21oi_1
XFILLER_21_784 VPWR VGND sg13g2_fill_1
XFILLER_0_633 VPWR VGND sg13g2_decap_8
X_6608__114 VPWR VGND net114 sg13g2_tiehi
XFILLER_43_342 VPWR VGND sg13g2_fill_1
XFILLER_15_1004 VPWR VGND sg13g2_decap_8
X_6615__107 VPWR VGND net107 sg13g2_tiehi
XFILLER_4_972 VPWR VGND sg13g2_decap_8
XFILLER_39_615 VPWR VGND sg13g2_fill_2
XFILLER_47_681 VPWR VGND sg13g2_fill_1
X_5901_ VGND VPWR _2561_ _2565_ _2567_ net424 sg13g2_a21oi_1
XFILLER_35_832 VPWR VGND sg13g2_fill_2
X_6881_ net323 VGND VPWR _0490_ u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[1\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_35_843 VPWR VGND sg13g2_fill_2
X_5832_ _2508_ _2507_ _2506_ VPWR VGND sg13g2_nand2b_1
X_5763_ VGND VPWR _2446_ _2449_ _0369_ _2450_ sg13g2_a21oi_1
X_4714_ _1579_ VPWR _1583_ VGND _1576_ _1581_ sg13g2_o21ai_1
X_5694_ VGND VPWR _2385_ _2390_ _2393_ _2389_ sg13g2_a21oi_1
XFILLER_30_581 VPWR VGND sg13g2_fill_2
X_6830__411 VPWR VGND net595 sg13g2_tiehi
X_4645_ VGND VPWR _1518_ _1520_ _1526_ _1525_ sg13g2_a21oi_1
Xhold700 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[7\] VPWR
+ VGND net1457 sg13g2_dlygate4sd3_1
Xhold711 _2339_ VPWR VGND net1468 sg13g2_dlygate4sd3_1
X_4576_ _1459_ VPWR _1468_ VGND net540 _0612_ sg13g2_o21ai_1
Xhold733 _0238_ VPWR VGND net1490 sg13g2_dlygate4sd3_1
X_6315_ _2895_ net758 net422 _2897_ VPWR VGND sg13g2_a21o_1
Xhold722 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[10\] VPWR VGND net1479
+ sg13g2_dlygate4sd3_1
X_3527_ VPWR _0597_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[8\]
+ VGND sg13g2_inv_1
Xhold755 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[9\] VPWR VGND net1512
+ sg13g2_dlygate4sd3_1
Xhold744 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[4\] VPWR VGND net1501
+ sg13g2_dlygate4sd3_1
Xhold766 _2694_ VPWR VGND net1523 sg13g2_dlygate4sd3_1
Xhold788 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[5\] VPWR VGND net1545
+ sg13g2_dlygate4sd3_1
Xhold777 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[8\].y_shr\[2\] VPWR
+ VGND net1534 sg13g2_dlygate4sd3_1
Xhold799 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[2\] VPWR VGND net1556
+ sg13g2_dlygate4sd3_1
X_6246_ _2853_ net510 net1099 VPWR VGND sg13g2_xnor2_1
X_6177_ _2796_ net1491 _2798_ VPWR VGND sg13g2_xor2_1
X_5128_ _1918_ _0566_ _1917_ VPWR VGND sg13g2_xnor2_1
X_6638__84 VPWR VGND net84 sg13g2_tiehi
X_6904__250 VPWR VGND net250 sg13g2_tiehi
X_5059_ VGND VPWR net1219 net395 _1871_ _1870_ sg13g2_a21oi_1
XFILLER_25_342 VPWR VGND sg13g2_fill_2
XFILLER_38_1026 VPWR VGND sg13g2_fill_2
XFILLER_21_570 VPWR VGND sg13g2_fill_2
XFILLER_4_213 VPWR VGND sg13g2_fill_2
XFILLER_5_758 VPWR VGND sg13g2_decap_8
XFILLER_1_931 VPWR VGND sg13g2_decap_8
XFILLER_49_924 VPWR VGND sg13g2_fill_1
Xhold60 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[1\] VPWR VGND net817
+ sg13g2_dlygate4sd3_1
Xhold71 u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[7\] VPWR VGND net828 sg13g2_dlygate4sd3_1
Xhold82 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[11\] VPWR VGND net839
+ sg13g2_dlygate4sd3_1
Xhold93 _0524_ VPWR VGND net850 sg13g2_dlygate4sd3_1
XFILLER_45_92 VPWR VGND sg13g2_fill_2
XFILLER_16_353 VPWR VGND sg13g2_fill_2
XFILLER_43_183 VPWR VGND sg13g2_fill_1
XFILLER_43_172 VPWR VGND sg13g2_fill_2
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk VPWR VGND sg13g2_buf_8
X_4430_ net433 _1345_ _1346_ _0139_ VPWR VGND sg13g2_nor3_1
X_6100_ _2731_ net1131 _2729_ VPWR VGND sg13g2_nand2_1
X_4361_ net436 _1288_ net1140 _0128_ VPWR VGND sg13g2_nor3_1
X_4292_ VPWR _1234_ net381 VGND sg13g2_inv_1
Xfanout509 net511 net509 VPWR VGND sg13g2_buf_2
X_6031_ _2671_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[3\] _2670_
+ VPWR VGND sg13g2_nand2_1
XFILLER_13_0 VPWR VGND sg13g2_fill_1
X_6635__87 VPWR VGND net87 sg13g2_tiehi
XFILLER_26_139 VPWR VGND sg13g2_fill_1
XFILLER_35_640 VPWR VGND sg13g2_fill_2
X_6864_ net357 VGND VPWR _0473_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[8\]
+ clknet_leaf_7_clk sg13g2_dfrbpq_2
X_5815_ _2491_ _2492_ _2493_ VPWR VGND sg13g2_nor2b_1
XFILLER_22_334 VPWR VGND sg13g2_fill_2
X_6795_ net630 VGND VPWR _0404_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[2\]
+ clknet_leaf_29_clk sg13g2_dfrbpq_1
X_5746_ VGND VPWR _2433_ _2435_ _0366_ _2436_ sg13g2_a21oi_1
X_5677_ _2377_ _2378_ _0355_ VPWR VGND sg13g2_nor2b_1
X_4628_ net1351 _1506_ _1511_ VPWR VGND sg13g2_nor2b_1
Xhold530 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[10\] VPWR
+ VGND net1287 sg13g2_dlygate4sd3_1
X_4559_ _1453_ VPWR _1454_ VGND net539 _0611_ sg13g2_o21ai_1
Xhold541 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[2\] VPWR
+ VGND net1298 sg13g2_dlygate4sd3_1
XFILLER_2_739 VPWR VGND sg13g2_decap_8
Xhold563 _2710_ VPWR VGND net1320 sg13g2_dlygate4sd3_1
Xhold552 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[10\] VPWR
+ VGND net1309 sg13g2_dlygate4sd3_1
Xhold585 _0222_ VPWR VGND net1342 sg13g2_dlygate4sd3_1
Xhold596 _0174_ VPWR VGND net1353 sg13g2_dlygate4sd3_1
Xhold574 _0445_ VPWR VGND net1331 sg13g2_dlygate4sd3_1
X_6229_ VGND VPWR _2835_ _2838_ _0446_ _2839_ sg13g2_a21oi_1
X_6605__117 VPWR VGND net117 sg13g2_tiehi
XFILLER_25_194 VPWR VGND sg13g2_fill_2
XFILLER_40_120 VPWR VGND sg13g2_fill_2
XFILLER_9_349 VPWR VGND sg13g2_fill_2
XFILLER_5_566 VPWR VGND sg13g2_fill_2
X_6820__421 VPWR VGND net605 sg13g2_tiehi
X_3930_ VGND VPWR _0533_ _0930_ _0932_ _0931_ sg13g2_a21oi_1
X_3861_ net441 VPWR _0891_ VGND net1019 _0888_ sg13g2_o21ai_1
XFILLER_16_194 VPWR VGND sg13g2_fill_1
X_6580_ net142 VGND VPWR net1294 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[5\]
+ clknet_leaf_34_clk sg13g2_dfrbpq_1
X_5600_ _2309_ VPWR _2312_ VGND _2306_ _2310_ sg13g2_o21ai_1
X_3792_ net882 u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[0\] _0839_ VPWR VGND sg13g2_xor2_1
X_5531_ VGND VPWR _2252_ _2253_ _0333_ _2254_ sg13g2_a21oi_1
XFILLER_9_883 VPWR VGND sg13g2_decap_8
X_5462_ VGND VPWR _2193_ _2197_ _0320_ _2198_ sg13g2_a21oi_1
X_5393_ net477 VPWR _2140_ VGND _2137_ _2139_ sg13g2_o21ai_1
X_4413_ VGND VPWR _1326_ _1331_ _1333_ net435 sg13g2_a21oi_1
X_4344_ _1276_ net502 _1275_ VPWR VGND sg13g2_nand2_1
X_6014_ VGND VPWR _2656_ _2655_ _0545_ sg13g2_or2_1
X_4275_ _1219_ _0585_ _1218_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_448 VPWR VGND sg13g2_fill_2
XFILLER_42_418 VPWR VGND sg13g2_fill_1
X_6916_ net266 VGND VPWR _0511_ u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[10\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_1
X_6847_ net578 VGND VPWR _0456_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[4\]
+ clknet_leaf_64_clk sg13g2_dfrbpq_2
XFILLER_11_805 VPWR VGND sg13g2_fill_2
XFILLER_23_676 VPWR VGND sg13g2_fill_1
X_6778_ net647 VGND VPWR _0387_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[11\]
+ clknet_leaf_58_clk sg13g2_dfrbpq_2
XFILLER_22_197 VPWR VGND sg13g2_fill_1
X_5729_ net491 VPWR _2424_ VGND _2422_ _2423_ sg13g2_o21ai_1
XFILLER_2_514 VPWR VGND sg13g2_fill_1
XFILLER_2_525 VPWR VGND sg13g2_fill_1
Xhold360 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[3\].y_shr\[8\] VPWR
+ VGND net1117 sg13g2_dlygate4sd3_1
Xhold371 _2470_ VPWR VGND net1128 sg13g2_dlygate4sd3_1
Xhold393 _1101_ VPWR VGND net1150 sg13g2_dlygate4sd3_1
Xhold382 _1287_ VPWR VGND net1139 sg13g2_dlygate4sd3_1
XFILLER_26_61 VPWR VGND sg13g2_fill_1
XFILLER_42_963 VPWR VGND sg13g2_fill_1
XFILLER_9_179 VPWR VGND sg13g2_fill_1
XFILLER_6_853 VPWR VGND sg13g2_decap_8
X_4060_ net1012 net548 net982 _1049_ VPWR VGND _1037_ sg13g2_nand4_1
XFILLER_37_702 VPWR VGND sg13g2_fill_1
XFILLER_18_982 VPWR VGND sg13g2_decap_8
X_4962_ _1789_ _1790_ _1788_ _1791_ VPWR VGND sg13g2_nand3_1
X_4893_ _1733_ net1251 net389 VPWR VGND sg13g2_nand2_1
X_3913_ net469 net800 _0043_ VPWR VGND sg13g2_and2_1
X_6701_ net724 VGND VPWR _0310_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[10\]
+ clknet_leaf_56_clk sg13g2_dfrbpq_2
X_6632_ net90 VGND VPWR net1397 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[5\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_1
X_3844_ net419 net951 _0878_ _0022_ VPWR VGND sg13g2_nor3_1
X_6563_ net159 VGND VPWR net1166 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[1\]
+ clknet_leaf_35_clk sg13g2_dfrbpq_2
X_3775_ net1019 u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[5\] net1023 _0822_ _0823_
+ VPWR VGND sg13g2_nor4_1
X_5514_ VGND VPWR _2241_ _2240_ _2238_ sg13g2_or2_1
X_6494_ net228 VGND VPWR _0103_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[1\]
+ clknet_leaf_45_clk sg13g2_dfrbpq_2
X_5445_ _2183_ _2178_ _2184_ VPWR VGND sg13g2_nor2b_1
X_5376_ VGND VPWR _0559_ _2118_ _2125_ net522 sg13g2_a21oi_1
X_4327_ net498 VPWR _1262_ VGND net770 _1261_ sg13g2_o21ai_1
X_4258_ _1204_ net1322 _1203_ VPWR VGND sg13g2_nand2_1
X_4189_ net534 _1137_ _1146_ VPWR VGND sg13g2_nor2_1
XFILLER_24_974 VPWR VGND sg13g2_decap_8
XFILLER_23_451 VPWR VGND sg13g2_fill_2
X_6810__431 VPWR VGND net615 sg13g2_tiehi
XFILLER_3_801 VPWR VGND sg13g2_decap_8
XFILLER_3_878 VPWR VGND sg13g2_decap_8
Xhold190 _1770_ VPWR VGND net947 sg13g2_dlygate4sd3_1
XFILLER_15_941 VPWR VGND sg13g2_decap_8
XFILLER_18_1024 VPWR VGND sg13g2_decap_4
X_3560_ net846 net446 _0525_ VPWR VGND sg13g2_and2_1
X_5230_ _1999_ net1538 _2003_ _2005_ VPWR VGND sg13g2_a21o_1
X_3491_ VPWR _0561_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[6\] VGND
+ sg13g2_inv_1
X_5161_ VGND VPWR _1944_ _1945_ _0271_ _1946_ sg13g2_a21oi_1
X_5092_ _1886_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[1\]
+ _1885_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_1017 VPWR VGND sg13g2_decap_8
XFILLER_25_1028 VPWR VGND sg13g2_fill_1
X_4112_ _1082_ _0582_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[6\]\[4\]
+ VPWR VGND sg13g2_nand2_1
X_4043_ _1036_ _0992_ _1034_ VPWR VGND sg13g2_nand2_1
X_5994_ _2637_ _2640_ _2635_ _2641_ VPWR VGND sg13g2_nand3_1
X_4945_ _1773_ VPWR _1776_ VGND _1769_ _1774_ sg13g2_o21ai_1
XFILLER_33_18 VPWR VGND sg13g2_fill_2
X_4876_ _1719_ net1447 _1717_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_933 VPWR VGND sg13g2_decap_8
X_6615_ net107 VGND VPWR _0224_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[11\]\[0\]
+ clknet_leaf_21_clk sg13g2_dfrbpq_1
X_3827_ _0866_ net552 _0867_ VPWR VGND _0865_ sg13g2_nand3b_1
X_6546_ net176 VGND VPWR net1478 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[9\]
+ clknet_leaf_38_clk sg13g2_dfrbpq_2
X_3758_ _0811_ _0806_ _0810_ VPWR VGND sg13g2_xnor2_1
X_3689_ VGND VPWR _0742_ _0741_ _0723_ sg13g2_or2_1
X_6477_ net245 VGND VPWR net1059 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[3\]
+ clknet_leaf_41_clk sg13g2_dfrbpq_1
X_5428_ VPWR _2169_ _2168_ VGND sg13g2_inv_1
XFILLER_0_815 VPWR VGND sg13g2_decap_8
X_5359_ VGND VPWR _0557_ _2094_ _2110_ net522 sg13g2_a21oi_1
XFILLER_15_259 VPWR VGND sg13g2_fill_1
XFILLER_12_900 VPWR VGND sg13g2_decap_8
XFILLER_8_937 VPWR VGND sg13g2_decap_8
XFILLER_12_977 VPWR VGND sg13g2_decap_8
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
XFILLER_48_70 VPWR VGND sg13g2_decap_8
XFILLER_48_81 VPWR VGND sg13g2_fill_2
X_6921__256 VPWR VGND net256 sg13g2_tiehi
X_4730_ _1597_ net1495 net400 VPWR VGND sg13g2_xnor2_1
X_4661_ _1524_ _1531_ _1518_ _1539_ VPWR VGND sg13g2_nand3_1
X_6400_ net563 VGND VPWR net897 net21 clknet_leaf_3_clk sg13g2_dfrbpq_2
X_3612_ _0658_ _0654_ _0665_ VPWR VGND sg13g2_xor2_1
X_4592_ VGND VPWR _1482_ _1481_ _1479_ sg13g2_or2_1
X_6331_ net763 net1007 _2898_ VPWR VGND sg13g2_and2_1
XFILLER_7_981 VPWR VGND sg13g2_decap_8
X_3543_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].z_sign _0613_ VPWR
+ VGND sg13g2_inv_4
X_3474_ VPWR _0544_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[10\]
+ VGND sg13g2_inv_1
X_6262_ net506 net1070 _2863_ _2864_ VPWR VGND sg13g2_nor3_1
X_5213_ _1986_ _1989_ _1990_ VPWR VGND sg13g2_nor2_1
X_6193_ _2812_ net1343 _2810_ VPWR VGND sg13g2_xnor2_1
X_5144_ net415 _0567_ _1932_ VPWR VGND sg13g2_nor2_1
X_5075_ net448 net3 _0249_ VPWR VGND sg13g2_and2_1
X_4026_ _1021_ net952 net377 VPWR VGND sg13g2_nand2_1
X_6800__441 VPWR VGND net625 sg13g2_tiehi
XFILLER_13_719 VPWR VGND sg13g2_fill_2
X_5977_ net467 net768 _0403_ VPWR VGND sg13g2_and2_1
X_4928_ net484 VPWR _1763_ VGND _1761_ _1762_ sg13g2_o21ai_1
X_4859_ net536 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[9\].y_shr\[0\]
+ _1704_ VPWR VGND sg13g2_nor2b_1
X_6529_ net193 VGND VPWR _0138_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[5\]
+ clknet_leaf_31_clk sg13g2_dfrbpq_1
XFILLER_0_689 VPWR VGND sg13g2_decap_8
XFILLER_18_95 VPWR VGND sg13g2_fill_1
XFILLER_12_774 VPWR VGND sg13g2_fill_2
XFILLER_4_951 VPWR VGND sg13g2_decap_8
X_5900_ _2561_ _2565_ _2566_ VPWR VGND sg13g2_nor2_1
XFILLER_34_321 VPWR VGND sg13g2_fill_2
X_6880_ net325 VGND VPWR _0489_ u_angle_cordic_12b_pmod.angle_cordic_12b.SINout\[0\]
+ clknet_leaf_22_clk sg13g2_dfrbpq_1
X_5831_ _2507_ _0578_ _2505_ VPWR VGND sg13g2_nand2_1
X_5762_ net472 VPWR _2450_ VGND _2446_ _2449_ sg13g2_o21ai_1
X_4713_ VGND VPWR _1576_ _1581_ _0187_ _1582_ sg13g2_a21oi_1
X_5693_ _2391_ _2392_ _0357_ VPWR VGND sg13g2_nor2b_1
X_4644_ _1525_ net1271 net393 VPWR VGND sg13g2_xnor2_1
Xhold701 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[7\] VPWR VGND net1458
+ sg13g2_dlygate4sd3_1
Xhold712 _0348_ VPWR VGND net1469 sg13g2_dlygate4sd3_1
X_4575_ _1462_ _1464_ _1467_ VPWR VGND sg13g2_nor2_1
X_3526_ _0596_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[5\] VPWR VGND
+ sg13g2_inv_2
Xhold734 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[8\] VPWR
+ VGND net1491 sg13g2_dlygate4sd3_1
Xhold745 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[4\].y_shr\[4\] VPWR
+ VGND net1502 sg13g2_dlygate4sd3_1
X_6314_ net758 _2895_ _2896_ VPWR VGND sg13g2_nor2_1
Xhold723 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[4\] VPWR
+ VGND net1480 sg13g2_dlygate4sd3_1
Xhold767 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[4\] VPWR VGND net1524
+ sg13g2_dlygate4sd3_1
X_6245_ _2850_ VPWR _2852_ VGND net510 _0563_ sg13g2_o21ai_1
Xhold756 _0117_ VPWR VGND net1513 sg13g2_dlygate4sd3_1
Xhold778 _1552_ VPWR VGND net1535 sg13g2_dlygate4sd3_1
Xhold789 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[3\] VPWR
+ VGND net1546 sg13g2_dlygate4sd3_1
X_6176_ net1491 _2796_ _2797_ VPWR VGND sg13g2_and2_1
X_5127_ net526 _1908_ _1917_ VPWR VGND sg13g2_nor2_1
XFILLER_29_126 VPWR VGND sg13g2_fill_1
X_5058_ net426 _1869_ net1220 _0244_ VPWR VGND sg13g2_nor3_1
XFILLER_26_822 VPWR VGND sg13g2_fill_2
X_4009_ _1007_ net954 net549 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_64_clk clknet_4_0_0_clk clknet_leaf_64_clk VPWR VGND sg13g2_buf_8
XFILLER_37_192 VPWR VGND sg13g2_fill_1
XFILLER_5_737 VPWR VGND sg13g2_decap_8
XFILLER_1_910 VPWR VGND sg13g2_decap_8
XFILLER_1_987 VPWR VGND sg13g2_decap_8
Xhold50 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[8\] VPWR VGND net807
+ sg13g2_dlygate4sd3_1
XFILLER_0_486 VPWR VGND sg13g2_fill_2
Xhold72 _0077_ VPWR VGND net829 sg13g2_dlygate4sd3_1
Xhold83 u_angle_cordic_12b_pmod.angle_cordic_12b.angle\[1\] VPWR VGND net840 sg13g2_dlygate4sd3_1
Xhold61 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[10\] VPWR VGND net818
+ sg13g2_dlygate4sd3_1
Xhold94 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.resetn VPWR VGND net851
+ sg13g2_dlygate4sd3_1
Xclkbuf_leaf_55_clk clknet_4_8_0_clk clknet_leaf_55_clk VPWR VGND sg13g2_buf_8
X_6621__101 VPWR VGND net101 sg13g2_tiehi
XFILLER_43_140 VPWR VGND sg13g2_fill_1
XFILLER_17_899 VPWR VGND sg13g2_decap_8
XFILLER_32_847 VPWR VGND sg13g2_fill_1
X_4360_ VGND VPWR _1283_ _1285_ _1289_ net1139 sg13g2_a21oi_1
X_4291_ VGND VPWR _1225_ _1233_ net1309 net531 sg13g2_a21oi_2
X_6030_ _2670_ _0620_ _2669_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_1014 VPWR VGND sg13g2_decap_8
XFILLER_20_2 VPWR VGND sg13g2_fill_1
XFILLER_26_107 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_46_clk clknet_4_11_0_clk clknet_leaf_46_clk VPWR VGND sg13g2_buf_8
X_6863_ net359 VGND VPWR _0472_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[7\]
+ clknet_leaf_2_clk sg13g2_dfrbpq_1
X_5814_ VGND VPWR _2492_ _2490_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[3\]
+ sg13g2_or2_1
XFILLER_23_858 VPWR VGND sg13g2_fill_2
X_6794_ net631 VGND VPWR _0403_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[1\]
+ clknet_leaf_28_clk sg13g2_dfrbpq_1
XFILLER_10_519 VPWR VGND sg13g2_fill_1
X_5745_ net468 VPWR _2436_ VGND _2433_ _2435_ sg13g2_o21ai_1
X_5676_ VGND VPWR _2371_ _2376_ _2378_ net431 sg13g2_a21oi_1
X_4627_ _1509_ net1350 _1510_ VPWR VGND sg13g2_xor2_1
Xhold520 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[2\] VPWR VGND net1277
+ sg13g2_dlygate4sd3_1
X_4558_ _0161_ net502 _1452_ _1453_ VPWR VGND sg13g2_and3_1
Xhold542 _0430_ VPWR VGND net1299 sg13g2_dlygate4sd3_1
XFILLER_2_718 VPWR VGND sg13g2_decap_8
Xhold553 _0107_ VPWR VGND net1310 sg13g2_dlygate4sd3_1
Xhold531 _0145_ VPWR VGND net1288 sg13g2_dlygate4sd3_1
Xhold575 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[7\]\[6\] VPWR VGND net1332
+ sg13g2_dlygate4sd3_1
X_3509_ VPWR _0579_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[6\] VGND
+ sg13g2_inv_1
Xhold564 _0422_ VPWR VGND net1321 sg13g2_dlygate4sd3_1
Xhold586 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[10\] VPWR
+ VGND net1343 sg13g2_dlygate4sd3_1
Xhold597 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[6\] VPWR VGND net1354
+ sg13g2_dlygate4sd3_1
X_4489_ _1397_ net1206 _1395_ VPWR VGND sg13g2_xnor2_1
X_6228_ net454 VPWR _2839_ VGND _2835_ _2838_ sg13g2_o21ai_1
X_6159_ _2782_ net1425 _2781_ VPWR VGND sg13g2_nand2b_1
Xclkbuf_leaf_37_clk clknet_4_15_0_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
XFILLER_26_630 VPWR VGND sg13g2_fill_2
XFILLER_12_1019 VPWR VGND sg13g2_decap_8
XFILLER_1_784 VPWR VGND sg13g2_decap_8
XFILLER_17_630 VPWR VGND sg13g2_fill_1
XFILLER_17_641 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_28_clk clknet_4_6_0_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
X_6894__545 VPWR VGND net729 sg13g2_tiehi
XFILLER_31_110 VPWR VGND sg13g2_fill_1
XFILLER_32_633 VPWR VGND sg13g2_fill_2
X_3860_ net1019 _0888_ _0890_ VPWR VGND sg13g2_and2_1
X_3791_ _0838_ u_angle_cordic_12b_pmod.u_vga_top.v_cnt\[9\] net835 VPWR VGND sg13g2_xnor2_1
XFILLER_9_862 VPWR VGND sg13g2_decap_8
X_5530_ net481 VPWR _2254_ VGND _2252_ _2253_ sg13g2_o21ai_1
X_5461_ net477 VPWR _2198_ VGND _2193_ _2197_ sg13g2_o21ai_1
X_4412_ _1326_ _1331_ _1332_ VPWR VGND sg13g2_nor2_1
X_5392_ _2133_ _2138_ _2139_ VPWR VGND sg13g2_nor2_1
X_4343_ VGND VPWR _1275_ _1274_ _1272_ sg13g2_or2_1
X_4274_ net531 _1210_ _1218_ VPWR VGND sg13g2_nor2_1
X_6013_ _2655_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[1\]
+ _2654_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_416 VPWR VGND sg13g2_fill_1
XFILLER_28_928 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_19_clk clknet_4_5_0_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
X_6915_ net268 VGND VPWR net848 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[9\]
+ clknet_leaf_15_clk sg13g2_dfrbpq_2
XFILLER_36_950 VPWR VGND sg13g2_fill_1
X_6631__91 VPWR VGND net91 sg13g2_tiehi
X_6846_ net579 VGND VPWR _0455_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[3\]
+ clknet_leaf_65_clk sg13g2_dfrbpq_2
X_6777_ net648 VGND VPWR net1424 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[3\]\[10\]
+ clknet_leaf_59_clk sg13g2_dfrbpq_2
X_3989_ _0990_ net940 net377 VPWR VGND sg13g2_nand2_1
X_5728_ _2423_ net1117 _2416_ VPWR VGND sg13g2_xnor2_1
X_5659_ VGND VPWR _2356_ _2361_ _2363_ net425 sg13g2_a21oi_1
X_6611__111 VPWR VGND net111 sg13g2_tiehi
Xhold361 _2423_ VPWR VGND net1118 sg13g2_dlygate4sd3_1
Xhold350 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt\[7\] VPWR VGND net1107
+ sg13g2_dlygate4sd3_1
Xhold372 _0374_ VPWR VGND net1129 sg13g2_dlygate4sd3_1
Xhold394 _1103_ VPWR VGND net1151 sg13g2_dlygate4sd3_1
Xhold383 _1289_ VPWR VGND net1140 sg13g2_dlygate4sd3_1
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk VPWR VGND sg13g2_buf_8
XFILLER_6_832 VPWR VGND sg13g2_decap_8
XFILLER_10_894 VPWR VGND sg13g2_decap_8
XFILLER_18_961 VPWR VGND sg13g2_decap_8
XFILLER_24_408 VPWR VGND sg13g2_fill_1
XFILLER_36_246 VPWR VGND sg13g2_fill_1
X_4961_ _1790_ net1112 net399 VPWR VGND sg13g2_xnor2_1
X_4892_ _1732_ _1730_ _1731_ VPWR VGND sg13g2_nand2_1
X_3912_ _0042_ net441 net792 net831 VPWR VGND sg13g2_and3_1
X_6700_ net739 VGND VPWR net1391 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[9\]
+ clknet_leaf_56_clk sg13g2_dfrbpq_2
X_6631_ net91 VGND VPWR _0240_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[4\]
+ clknet_leaf_20_clk sg13g2_dfrbpq_1
X_3843_ net950 _0876_ _0878_ VPWR VGND sg13g2_and2_1
X_6562_ net160 VGND VPWR _0171_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[0\]
+ clknet_leaf_37_clk sg13g2_dfrbpq_2
X_3774_ u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[10\] u_angle_cordic_12b_pmod.u_vga_top.h_cnt\[9\]
+ _0540_ _0822_ VPWR VGND sg13g2_or3_1
X_5513_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[4\] net523 _2240_
+ VPWR VGND sg13g2_xor2_1
X_6493_ net229 VGND VPWR _0102_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[7\].y_shr\[0\]
+ clknet_leaf_45_clk sg13g2_dfrbpq_2
X_5444_ _2180_ net1317 _2183_ VPWR VGND sg13g2_xor2_1
Xclkbuf_leaf_8_clk clknet_4_3_0_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_5375_ _2121_ VPWR _2124_ VGND _2117_ _2122_ sg13g2_o21ai_1
X_4326_ _1261_ net542 net817 VPWR VGND sg13g2_xnor2_1
X_4257_ _1202_ net1576 _1203_ VPWR VGND sg13g2_xor2_1
X_4188_ _1141_ _1136_ _1140_ _1145_ VPWR VGND sg13g2_a21o_2
XFILLER_24_953 VPWR VGND sg13g2_decap_8
X_6829_ net596 VGND VPWR net1345 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[2\].y_shr\[9\]
+ clknet_leaf_8_clk sg13g2_dfrbpq_2
XFILLER_3_857 VPWR VGND sg13g2_decap_8
Xhold180 _0879_ VPWR VGND net937 sg13g2_dlygate4sd3_1
Xhold191 u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp\[4\] VPWR VGND
+ net948 sg13g2_dlygate4sd3_1
XFILLER_15_920 VPWR VGND sg13g2_decap_8
XFILLER_33_216 VPWR VGND sg13g2_fill_1
XFILLER_18_1003 VPWR VGND sg13g2_decap_8
XFILLER_15_997 VPWR VGND sg13g2_decap_8
X_3490_ VPWR _0560_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[4\]\[8\] VGND
+ sg13g2_inv_1
X_5160_ net492 VPWR _1946_ VGND _1944_ _1945_ sg13g2_o21ai_1
X_5091_ _1885_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[5\].y_shr\[0\]
+ net526 VPWR VGND sg13g2_nand2b_1
X_4111_ VGND VPWR _1077_ net1058 _0086_ _1081_ sg13g2_a21oi_1
X_6861__363 VPWR VGND net363 sg13g2_tiehi
X_4042_ _1035_ _1033_ _1028_ _1032_ _0939_ VPWR VGND sg13g2_a22oi_1
XFILLER_37_500 VPWR VGND sg13g2_fill_1
XFILLER_37_566 VPWR VGND sg13g2_fill_2
X_5993_ net1325 net513 _2640_ VPWR VGND sg13g2_xor2_1
X_4944_ VGND VPWR _1769_ _1774_ _0225_ _1775_ sg13g2_a21oi_1
X_6601__121 VPWR VGND net121 sg13g2_tiehi
XFILLER_33_750 VPWR VGND sg13g2_fill_1
X_4875_ _1717_ net1447 _1718_ VPWR VGND sg13g2_nor2b_1
X_6614_ net108 VGND VPWR net1216 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[10\]\[12\]
+ clknet_leaf_25_clk sg13g2_dfrbpq_2
X_3826_ _0864_ VPWR _0866_ VGND _0812_ _0816_ sg13g2_o21ai_1
XFILLER_21_989 VPWR VGND sg13g2_decap_8
X_6545_ net177 VGND VPWR _0154_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[8\]
+ clknet_leaf_37_clk sg13g2_dfrbpq_2
X_3757_ _0809_ VPWR _0810_ VGND _0772_ _0808_ sg13g2_o21ai_1
X_6476_ net246 VGND VPWR _0085_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[7\]\[2\]
+ clknet_leaf_41_clk sg13g2_dfrbpq_1
X_3688_ VPWR VGND _0737_ _0740_ _0735_ _0717_ _0741_ _0722_ sg13g2_a221oi_1
X_5427_ _2166_ net1367 _2168_ VPWR VGND sg13g2_xor2_1
X_5358_ _2106_ VPWR _2109_ VGND _2103_ _2107_ sg13g2_o21ai_1
X_4309_ _1234_ VPWR _1248_ VGND u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[8\]
+ net1512 sg13g2_o21ai_1
X_5289_ _2052_ net496 _2051_ VPWR VGND sg13g2_nand2_1
XFILLER_12_956 VPWR VGND sg13g2_decap_8
XFILLER_8_916 VPWR VGND sg13g2_decap_8
XFILLER_7_415 VPWR VGND sg13g2_fill_1
XFILLER_48_1007 VPWR VGND sg13g2_decap_8
Xfanout490 net491 net490 VPWR VGND sg13g2_buf_8
X_6409__362 VPWR VGND net362 sg13g2_tiehi
X_4660_ VGND VPWR _0610_ _1523_ _1538_ _1532_ sg13g2_a21oi_1
X_3611_ VPWR _0664_ _0663_ VGND sg13g2_inv_1
XFILLER_7_960 VPWR VGND sg13g2_decap_8
X_6330_ net763 net374 _0501_ VPWR VGND sg13g2_nor2_1
X_4591_ net1086 net540 _1481_ VPWR VGND sg13g2_xor2_1
X_3542_ VPWR _0612_ net1153 VGND sg13g2_inv_1
X_3473_ _0543_ net1041 VPWR VGND sg13g2_inv_2
X_6261_ net967 net555 _2863_ VPWR VGND sg13g2_nor2_1
X_5212_ net439 _1988_ _1989_ _0279_ VPWR VGND sg13g2_nor3_1
X_6192_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[10\] _2810_
+ _2811_ VPWR VGND sg13g2_and2_1
XFILLER_9_1023 VPWR VGND sg13g2_decap_4
X_5143_ _1925_ net1162 _1929_ _1931_ VPWR VGND sg13g2_a21o_1
X_5074_ net448 net2 _0248_ VPWR VGND sg13g2_and2_1
X_4025_ _1015_ VPWR _0061_ VGND net372 _1020_ sg13g2_o21ai_1
X_5976_ net467 net791 _0402_ VPWR VGND sg13g2_and2_1
X_4927_ _1752_ _1758_ _1762_ VPWR VGND sg13g2_and2_1
XFILLER_21_742 VPWR VGND sg13g2_fill_2
X_4858_ net999 _1702_ _0211_ VPWR VGND sg13g2_nor2b_1
X_3809_ net553 net892 _0852_ VPWR VGND sg13g2_nor2_1
X_4789_ VGND VPWR _0613_ _1645_ _1646_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[9\]\[11\]
+ sg13g2_a21oi_1
XFILLER_5_919 VPWR VGND sg13g2_decap_8
X_6528_ net194 VGND VPWR net1376 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[8\]\[4\]
+ clknet_leaf_41_clk sg13g2_dfrbpq_2
X_6459_ net275 VGND VPWR _0068_ u_angle_cordic_12b_pmod.waveform_sel_reg\[0\] clknet_leaf_16_clk
+ sg13g2_dfrbpq_2
XFILLER_0_668 VPWR VGND sg13g2_decap_8
XFILLER_18_41 VPWR VGND sg13g2_fill_2
XFILLER_29_897 VPWR VGND sg13g2_fill_2
XFILLER_16_536 VPWR VGND sg13g2_fill_2
XFILLER_16_547 VPWR VGND sg13g2_fill_1
XFILLER_4_930 VPWR VGND sg13g2_decap_8
XFILLER_3_451 VPWR VGND sg13g2_fill_1
XFILLER_39_617 VPWR VGND sg13g2_fill_1
X_6647__75 VPWR VGND net75 sg13g2_tiehi
XFILLER_38_116 VPWR VGND sg13g2_fill_2
X_5830_ _0578_ _2505_ _2506_ VPWR VGND sg13g2_nor2_1
XFILLER_22_539 VPWR VGND sg13g2_fill_1
X_5761_ _2449_ net518 net1084 VPWR VGND sg13g2_xnor2_1
X_4712_ net488 VPWR _1582_ VGND _1576_ _1581_ sg13g2_o21ai_1
X_5692_ VGND VPWR _2385_ _2390_ _2392_ net431 sg13g2_a21oi_1
X_4643_ _1524_ net1550 net393 VPWR VGND sg13g2_nand2_1
Xhold702 _1609_ VPWR VGND net1459 sg13g2_dlygate4sd3_1
X_4574_ net436 _1465_ _1466_ _0164_ VPWR VGND sg13g2_nor3_1
Xhold713 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[9\]\[2\] VPWR VGND net1470
+ sg13g2_dlygate4sd3_1
Xhold724 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[4\] VPWR VGND net1481
+ sg13g2_dlygate4sd3_1
X_6313_ _2895_ net506 net815 VPWR VGND sg13g2_xnor2_1
X_3525_ _0595_ net1519 VPWR VGND sg13g2_inv_2
Xhold735 _0436_ VPWR VGND net1492 sg13g2_dlygate4sd3_1
Xhold746 _0322_ VPWR VGND net1503 sg13g2_dlygate4sd3_1
Xhold779 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[7\] VPWR
+ VGND net1536 sg13g2_dlygate4sd3_1
X_6244_ VGND VPWR net1072 _2849_ _0449_ _2851_ sg13g2_a21oi_1
Xhold768 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[7\]\[2\] VPWR VGND net1525
+ sg13g2_dlygate4sd3_1
Xhold757 u_angle_cordic_12b_pmod.waveform_sel_reg\[1\] VPWR VGND net1514 sg13g2_dlygate4sd3_1
X_6175_ _2796_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[10\] _2794_
+ VPWR VGND sg13g2_xnor2_1
X_5126_ _1916_ _1910_ _1915_ VPWR VGND sg13g2_nand2_1
X_5057_ VGND VPWR _1865_ _1867_ _1870_ _1868_ sg13g2_a21oi_1
X_4008_ net954 net550 _1006_ VPWR VGND sg13g2_nor2_1
XFILLER_38_1028 VPWR VGND sg13g2_fill_1
X_5959_ _2617_ net1530 _2616_ VPWR VGND sg13g2_nand2_1
XFILLER_5_716 VPWR VGND sg13g2_decap_8
XFILLER_4_215 VPWR VGND sg13g2_fill_1
X_6911__278 VPWR VGND net278 sg13g2_tiehi
XFILLER_1_966 VPWR VGND sg13g2_decap_8
Xhold40 _0496_ VPWR VGND net797 sg13g2_dlygate4sd3_1
Xhold51 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[11\]\[5\] VPWR VGND net808
+ sg13g2_dlygate4sd3_1
XFILLER_21_1010 VPWR VGND sg13g2_decap_8
Xhold62 _0132_ VPWR VGND net819 sg13g2_dlygate4sd3_1
Xhold73 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[5\]\[1\] VPWR VGND net830
+ sg13g2_dlygate4sd3_1
XFILLER_17_812 VPWR VGND sg13g2_fill_1
Xhold84 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[2\]\[6\] VPWR VGND net841
+ sg13g2_dlygate4sd3_1
X_6644__78 VPWR VGND net78 sg13g2_tiehi
Xhold95 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[4\]\[0\] VPWR VGND net852
+ sg13g2_dlygate4sd3_1
XFILLER_12_550 VPWR VGND sg13g2_fill_1
X_4290_ VGND VPWR _1223_ _1229_ _1232_ _1227_ sg13g2_a21oi_1
X_6862_ net361 VGND VPWR _0471_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[6\]
+ clknet_leaf_63_clk sg13g2_dfrbpq_2
X_5813_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[2\]\[3\] _2490_ _2491_
+ VPWR VGND sg13g2_and2_1
X_6793_ net632 VGND VPWR _0402_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[3\]\[0\]
+ clknet_leaf_28_clk sg13g2_dfrbpq_1
X_5744_ net1280 net517 _2435_ VPWR VGND sg13g2_xor2_1
X_5675_ _2371_ _2376_ _2377_ VPWR VGND sg13g2_nor2_1
XFILLER_30_391 VPWR VGND sg13g2_fill_1
X_4626_ _1509_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[11\] _1508_
+ VPWR VGND sg13g2_xnor2_1
Xhold510 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z\[1\]\[7\] VPWR VGND net1267
+ sg13g2_dlygate4sd3_1
X_4557_ _1449_ _1447_ _1451_ _1453_ VPWR VGND sg13g2_a21o_1
Xhold554 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[8\]\[3\] VPWR VGND net1311
+ sg13g2_dlygate4sd3_1
Xhold532 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[5\]\[9\] VPWR VGND net1289
+ sg13g2_dlygate4sd3_1
Xhold521 _1198_ VPWR VGND net1278 sg13g2_dlygate4sd3_1
Xhold543 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[6\].y_shr\[4\] VPWR
+ VGND net1300 sg13g2_dlygate4sd3_1
Xhold576 _0153_ VPWR VGND net1333 sg13g2_dlygate4sd3_1
X_3508_ VPWR _0578_ net1553 VGND sg13g2_inv_1
Xhold587 _2812_ VPWR VGND net1344 sg13g2_dlygate4sd3_1
Xhold565 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[6\]\[3\] VPWR VGND net1322
+ sg13g2_dlygate4sd3_1
X_4488_ _1396_ net1206 _1395_ VPWR VGND sg13g2_nand2_1
Xhold598 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y\[6\]\[2\] VPWR VGND net1355
+ sg13g2_dlygate4sd3_1
X_6227_ _2838_ _2837_ _2836_ VPWR VGND sg13g2_nand2b_1
X_6158_ _2779_ u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x\[1\]\[8\] _2781_
+ VPWR VGND sg13g2_xor2_1
X_5109_ _1901_ _0565_ _1900_ VPWR VGND sg13g2_xnor2_1
X_6089_ _2722_ _2714_ _2717_ _2721_ VPWR VGND sg13g2_and3_1
X_6464__267 VPWR VGND net267 sg13g2_tiehi
XFILLER_26_686 VPWR VGND sg13g2_fill_1
XFILLER_40_122 VPWR VGND sg13g2_fill_1
XFILLER_5_502 VPWR VGND sg13g2_fill_1
XFILLER_5_568 VPWR VGND sg13g2_fill_1
XFILLER_31_96 VPWR VGND sg13g2_fill_1
XFILLER_1_763 VPWR VGND sg13g2_decap_8
XFILLER_0_273 VPWR VGND sg13g2_fill_2
XFILLER_44_461 VPWR VGND sg13g2_fill_2
XFILLER_13_881 VPWR VGND sg13g2_decap_8
X_3790_ VPWR VGND _0534_ _0834_ net889 net1003 _0837_ _0550_ sg13g2_a221oi_1
XFILLER_20_829 VPWR VGND sg13g2_fill_2
XFILLER_9_841 VPWR VGND sg13g2_decap_8
XFILLER_8_373 VPWR VGND sg13g2_fill_2
X_5460_ _2197_ net1388 _2195_ VPWR VGND sg13g2_xnor2_1
X_4411_ _1329_ net1374 _1331_ VPWR VGND sg13g2_xor2_1
X_5391_ VPWR VGND net1390 _2127_ _2132_ _2124_ _2138_ _2128_ sg13g2_a221oi_1
X_4342_ net1080 net541 _1274_ VPWR VGND sg13g2_xor2_1
X_4273_ VGND VPWR _1207_ _1213_ _1217_ _1212_ sg13g2_a21oi_1
XFILLER_28_1027 VPWR VGND sg13g2_fill_2
X_6012_ net507 u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz\[1\].y_shr\[0\]
+ _2654_ VPWR VGND sg13g2_nor2b_1
.ends

