module heichips25_CORDIC (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire hsync_sig;
 wire pwm_data;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle[11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle[3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle[4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle[5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle[6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle[7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle[8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle[9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[12] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[13] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[14] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[15] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[16] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[17] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt_sum[5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[12] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.resetn ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp[11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.up ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.x_start[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[0][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][12] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][12] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][12] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][12] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][12] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][12] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][12] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][12] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][12] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][12] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[0].y_shr[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[0].y_shr[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[0].y_shr[11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[0].z_sign ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].z_sign ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].z_sign ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].z_sign ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].z_sign ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].z_sign ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].z_sign ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].z_sign ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].z_sign ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].z_sign ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].z_sign ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][11] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[2][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[2][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[3][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[3][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[3][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[4][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[4][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[4][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[4][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][9] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][0] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][10] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][1] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][2] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][3] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][4] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][5] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][6] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][7] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][8] ;
 wire \u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][9] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.clk_div_cnt[0] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.clk_div_cnt[1] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.h_cnt[0] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.h_cnt[10] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.h_cnt[1] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.h_cnt[2] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.h_cnt[3] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.h_cnt[4] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.h_cnt[5] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.h_cnt[6] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.h_cnt[7] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.h_cnt[8] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.h_cnt[9] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.pixel_clk_en ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_cnt[0] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_cnt[10] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_cnt[1] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_cnt[2] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_cnt[3] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_cnt[4] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_cnt[5] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_cnt[6] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_cnt[7] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_cnt[8] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_cnt[9] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_pos[0] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_pos[10] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_pos[1] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_pos[2] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_pos[3] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_pos[4] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_pos[5] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_pos[6] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_pos[7] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_pos[8] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.v_pos[9] ;
 wire \u_angle_cordic_12b_pmod.u_vga_top.vsync ;
 wire \u_angle_cordic_12b_pmod.waveform_sel_reg[0] ;
 wire \u_angle_cordic_12b_pmod.waveform_sel_reg[1] ;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire clknet_leaf_0_clk;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net17;
 wire net18;
 wire net19;
 wire net39;
 wire net20;
 wire net21;
 wire net22;
 wire net40;
 wire net23;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net24;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;

 sg13g2_inv_1 _3461_ (.Y(_0531_),
    .A(net856));
 sg13g2_inv_1 _3462_ (.Y(_0532_),
    .A(net803));
 sg13g2_inv_1 _3463_ (.Y(_0533_),
    .A(net885));
 sg13g2_inv_1 _3464_ (.Y(_0534_),
    .A(net914));
 sg13g2_inv_1 _3465_ (.Y(_0535_),
    .A(net978));
 sg13g2_inv_1 _3466_ (.Y(_0536_),
    .A(net920));
 sg13g2_inv_1 _3467_ (.Y(_0537_),
    .A(net1024));
 sg13g2_inv_1 _3468_ (.Y(_0538_),
    .A(net983));
 sg13g2_inv_2 _3469_ (.Y(_0539_),
    .A(net554));
 sg13g2_inv_1 _3470_ (.Y(_0540_),
    .A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[8] ));
 sg13g2_inv_1 _3471_ (.Y(_0541_),
    .A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[7] ));
 sg13g2_inv_1 _3472_ (.Y(_0542_),
    .A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[6] ));
 sg13g2_inv_2 _3473_ (.Y(_0543_),
    .A(net1041));
 sg13g2_inv_1 _3474_ (.Y(_0544_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][10] ));
 sg13g2_inv_1 _3475_ (.Y(_0545_),
    .A(net965));
 sg13g2_inv_1 _3476_ (.Y(_0546_),
    .A(net459));
 sg13g2_inv_1 _3477_ (.Y(_0547_),
    .A(net1107));
 sg13g2_inv_1 _3478_ (.Y(_0548_),
    .A(net892));
 sg13g2_inv_1 _3479_ (.Y(_0549_),
    .A(net909));
 sg13g2_inv_1 _3480_ (.Y(_0550_),
    .A(net944));
 sg13g2_inv_1 _3481_ (.Y(_0551_),
    .A(net929));
 sg13g2_inv_1 _3482_ (.Y(_0552_),
    .A(net889));
 sg13g2_inv_2 _3483_ (.Y(_0553_),
    .A(net523));
 sg13g2_inv_1 _3484_ (.Y(_0554_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][1] ));
 sg13g2_inv_2 _3485_ (.Y(_0555_),
    .A(net1566));
 sg13g2_inv_1 _3486_ (.Y(_0556_),
    .A(net1517));
 sg13g2_inv_2 _3487_ (.Y(_0557_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[5] ));
 sg13g2_inv_1 _3488_ (.Y(_0558_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][6] ));
 sg13g2_inv_2 _3489_ (.Y(_0559_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[7] ));
 sg13g2_inv_1 _3490_ (.Y(_0560_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][8] ));
 sg13g2_inv_1 _3491_ (.Y(_0561_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][6] ));
 sg13g2_inv_1 _3492_ (.Y(_0562_),
    .A(net509));
 sg13g2_inv_1 _3493_ (.Y(_0563_),
    .A(net1392));
 sg13g2_inv_1 _3494_ (.Y(_0564_),
    .A(net529));
 sg13g2_inv_2 _3495_ (.Y(_0565_),
    .A(net1181));
 sg13g2_inv_1 _3496_ (.Y(_0566_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[5] ));
 sg13g2_inv_2 _3497_ (.Y(_0567_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[10] ));
 sg13g2_inv_2 _3498_ (.Y(_0568_),
    .A(net1410));
 sg13g2_inv_1 _3499_ (.Y(_0569_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][8] ));
 sg13g2_inv_1 _3500_ (.Y(_0570_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][9] ));
 sg13g2_inv_2 _3501_ (.Y(_0571_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][10] ));
 sg13g2_inv_1 _3502_ (.Y(_0572_),
    .A(net1259));
 sg13g2_inv_1 _3503_ (.Y(_0573_),
    .A(net512));
 sg13g2_inv_1 _3504_ (.Y(_0574_),
    .A(net1427));
 sg13g2_inv_1 _3505_ (.Y(_0575_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[2] ));
 sg13g2_inv_1 _3506_ (.Y(_0576_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][4] ));
 sg13g2_inv_1 _3507_ (.Y(_0577_),
    .A(net1554));
 sg13g2_inv_1 _3508_ (.Y(_0578_),
    .A(net1553));
 sg13g2_inv_1 _3509_ (.Y(_0579_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][6] ));
 sg13g2_inv_1 _3510_ (.Y(_0580_),
    .A(net1562));
 sg13g2_inv_1 _3511_ (.Y(_0581_),
    .A(net1531));
 sg13g2_inv_4 _3512_ (.A(net531),
    .Y(_0582_));
 sg13g2_inv_1 _3513_ (.Y(_0583_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][1] ));
 sg13g2_inv_1 _3514_ (.Y(_0584_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[2] ));
 sg13g2_inv_1 _3515_ (.Y(_0585_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[5] ));
 sg13g2_inv_1 _3516_ (.Y(_0586_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][8] ));
 sg13g2_inv_1 _3517_ (.Y(_0587_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][11] ));
 sg13g2_inv_1 _3518_ (.Y(_0588_),
    .A(net1154));
 sg13g2_inv_1 _3519_ (.Y(_0589_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][6] ));
 sg13g2_inv_1 _3520_ (.Y(_0590_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][8] ));
 sg13g2_inv_1 _3521_ (.Y(_0591_),
    .A(net1115));
 sg13g2_inv_2 _3522_ (.Y(_0592_),
    .A(net519));
 sg13g2_inv_1 _3523_ (.Y(_0593_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][1] ));
 sg13g2_inv_1 _3524_ (.Y(_0594_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[2] ));
 sg13g2_inv_2 _3525_ (.Y(_0595_),
    .A(net1519));
 sg13g2_inv_2 _3526_ (.Y(_0596_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][5] ));
 sg13g2_inv_1 _3527_ (.Y(_0597_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[8] ));
 sg13g2_inv_2 _3528_ (.Y(_0598_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[10] ));
 sg13g2_inv_1 _3529_ (.Y(_0599_),
    .A(net1482));
 sg13g2_inv_1 _3530_ (.Y(_0600_),
    .A(net541));
 sg13g2_inv_1 _3531_ (.Y(_0601_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[3] ));
 sg13g2_inv_1 _3532_ (.Y(_0602_),
    .A(net1441));
 sg13g2_inv_1 _3533_ (.Y(_0603_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][10] ));
 sg13g2_inv_2 _3534_ (.Y(_0604_),
    .A(net1525));
 sg13g2_inv_1 _3535_ (.Y(_0605_),
    .A(net506));
 sg13g2_inv_1 _3536_ (.Y(_0606_),
    .A(net1120));
 sg13g2_inv_1 _3537_ (.Y(_0607_),
    .A(net1110));
 sg13g2_inv_2 _3538_ (.Y(_0608_),
    .A(net540));
 sg13g2_inv_1 _3539_ (.Y(_0609_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[2] ));
 sg13g2_inv_1 _3540_ (.Y(_0610_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][7] ));
 sg13g2_inv_1 _3541_ (.Y(_0611_),
    .A(net1272));
 sg13g2_inv_1 _3542_ (.Y(_0612_),
    .A(net1153));
 sg13g2_inv_4 _3543_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].z_sign ),
    .Y(_0613_));
 sg13g2_inv_1 _3544_ (.Y(_0614_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][1] ));
 sg13g2_inv_1 _3545_ (.Y(_0615_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[2] ));
 sg13g2_inv_1 _3546_ (.Y(_0616_),
    .A(net1556));
 sg13g2_inv_1 _3547_ (.Y(_0617_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].z_sign ));
 sg13g2_inv_1 _3548_ (.Y(_0618_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][4] ));
 sg13g2_inv_1 _3549_ (.Y(_0619_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][3] ));
 sg13g2_inv_2 _3550_ (.Y(_0620_),
    .A(net1546));
 sg13g2_inv_1 _3551_ (.Y(_0621_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][7] ));
 sg13g2_inv_1 _3552_ (.Y(_0622_),
    .A(net1536));
 sg13g2_inv_1 _3553_ (.Y(_0623_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][9] ));
 sg13g2_inv_1 _3554_ (.Y(_0624_),
    .A(net1130));
 sg13g2_inv_1 _3555_ (.Y(_0625_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[10] ));
 sg13g2_and2_1 _3556_ (.A(net879),
    .B(net451),
    .X(_0519_));
 sg13g2_and2_1 _3557_ (.A(net840),
    .B(net450),
    .X(_0522_));
 sg13g2_and2_1 _3558_ (.A(net919),
    .B(net450),
    .X(_0523_));
 sg13g2_and2_1 _3559_ (.A(net849),
    .B(net451),
    .X(_0524_));
 sg13g2_and2_1 _3560_ (.A(net846),
    .B(net446),
    .X(_0525_));
 sg13g2_and2_1 _3561_ (.A(net824),
    .B(net445),
    .X(_0526_));
 sg13g2_nor2_1 _3562_ (.A(_0531_),
    .B(net422),
    .Y(_0527_));
 sg13g2_and2_1 _3563_ (.A(net828),
    .B(net445),
    .X(_0528_));
 sg13g2_and2_1 _3564_ (.A(net821),
    .B(net445),
    .X(_0529_));
 sg13g2_and2_1 _3565_ (.A(net865),
    .B(net444),
    .X(_0530_));
 sg13g2_and2_1 _3566_ (.A(net878),
    .B(net442),
    .X(_0520_));
 sg13g2_nand3_1 _3567_ (.B(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[5] ),
    .C(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[4] ),
    .A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[6] ),
    .Y(_0626_));
 sg13g2_nand2_1 _3568_ (.Y(_0627_),
    .A(_0538_),
    .B(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[9] ));
 sg13g2_nor3_1 _3569_ (.A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[6] ),
    .B(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[5] ),
    .C(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[4] ),
    .Y(_0628_));
 sg13g2_nor4_1 _3570_ (.A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[8] ),
    .B(_0541_),
    .C(_0627_),
    .D(_0628_),
    .Y(_0629_));
 sg13g2_nand2_1 _3571_ (.Y(hsync_sig),
    .A(_0626_),
    .B(_0629_));
 sg13g2_and4_1 _3572_ (.A(net914),
    .B(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[7] ),
    .C(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[6] ),
    .D(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[5] ),
    .X(_0630_));
 sg13g2_nor4_1 _3573_ (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[10] ),
    .B(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[9] ),
    .C(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[4] ),
    .D(_0535_),
    .Y(_0631_));
 sg13g2_nand2_1 _3574_ (.Y(_0632_),
    .A(net978),
    .B(net920));
 sg13g2_nand4_1 _3575_ (.B(_0630_),
    .C(_0631_),
    .A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[1] ),
    .Y(\u_angle_cordic_12b_pmod.u_vga_top.vsync ),
    .D(_0632_));
 sg13g2_nand2_1 _3576_ (.Y(_0633_),
    .A(net442),
    .B(net822));
 sg13g2_nand2b_1 _3577_ (.Y(_0634_),
    .B(net878),
    .A_N(net859));
 sg13g2_nor2_1 _3578_ (.A(_0633_),
    .B(_0634_),
    .Y(_0000_));
 sg13g2_nand2b_1 _3579_ (.Y(_0635_),
    .B(net859),
    .A_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[11] ));
 sg13g2_nor2_1 _3580_ (.A(_0633_),
    .B(net860),
    .Y(_0001_));
 sg13g2_a21oi_1 _3581_ (.A1(_0634_),
    .A2(net860),
    .Y(_0002_),
    .B1(_0633_));
 sg13g2_and4_1 _3582_ (.A(net442),
    .B(net822),
    .C(_0634_),
    .D(_0635_),
    .X(_0003_));
 sg13g2_mux4_1 _3583_ (.S0(\u_angle_cordic_12b_pmod.waveform_sel_reg[0] ),
    .A0(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[11] ),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[11] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[11] ),
    .A3(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp[11] ),
    .S1(net1514),
    .X(_0636_));
 sg13g2_mux4_1 _3584_ (.S0(net546),
    .A0(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[1] ),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[1] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[1] ),
    .A3(net535),
    .S1(net544),
    .X(_0637_));
 sg13g2_mux4_1 _3585_ (.S0(net546),
    .A0(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[2] ),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[2] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[2] ),
    .A3(net535),
    .S1(net544),
    .X(_0638_));
 sg13g2_mux4_1 _3586_ (.S0(net547),
    .A0(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[0] ),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[0] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[0] ),
    .A3(net535),
    .S1(net545),
    .X(_0639_));
 sg13g2_mux4_1 _3587_ (.S0(net546),
    .A0(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[3] ),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[3] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[3] ),
    .A3(net535),
    .S1(net544),
    .X(_0640_));
 sg13g2_mux4_1 _3588_ (.S0(net546),
    .A0(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[6] ),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[6] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[6] ),
    .A3(net535),
    .S1(net544),
    .X(_0641_));
 sg13g2_mux4_1 _3589_ (.S0(net546),
    .A0(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[7] ),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[7] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[7] ),
    .A3(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp[0] ),
    .S1(net544),
    .X(_0642_));
 sg13g2_mux4_1 _3590_ (.S0(net546),
    .A0(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[5] ),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[5] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[5] ),
    .A3(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp[11] ),
    .S1(net544),
    .X(_0643_));
 sg13g2_mux4_1 _3591_ (.S0(net547),
    .A0(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[4] ),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[4] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[4] ),
    .A3(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp[11] ),
    .S1(net545),
    .X(_0644_));
 sg13g2_nor2_1 _3592_ (.A(net407),
    .B(net406),
    .Y(_0645_));
 sg13g2_mux4_1 _3593_ (.S0(net546),
    .A0(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[9] ),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[9] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[9] ),
    .A3(net535),
    .S1(net544),
    .X(_0646_));
 sg13g2_mux4_1 _3594_ (.S0(net546),
    .A0(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[8] ),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[8] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[8] ),
    .A3(net535),
    .S1(net544),
    .X(_0647_));
 sg13g2_or2_1 _3595_ (.X(_0648_),
    .B(_0639_),
    .A(_0637_));
 sg13g2_nor4_1 _3596_ (.A(_0638_),
    .B(_0640_),
    .C(net407),
    .D(net406),
    .Y(_0649_));
 sg13g2_nor4_1 _3597_ (.A(_0641_),
    .B(net408),
    .C(net404),
    .D(net403),
    .Y(_0650_));
 sg13g2_nand3b_1 _3598_ (.B(_0649_),
    .C(_0650_),
    .Y(_0651_),
    .A_N(_0648_));
 sg13g2_nand2_1 _3599_ (.Y(_0652_),
    .A(_0636_),
    .B(_0651_));
 sg13g2_xor2_1 _3600_ (.B(net408),
    .A(net409),
    .X(_0653_));
 sg13g2_nand2_1 _3601_ (.Y(_0654_),
    .A(_0637_),
    .B(_0653_));
 sg13g2_and2_1 _3602_ (.A(net408),
    .B(net403),
    .X(_0655_));
 sg13g2_xor2_1 _3603_ (.B(net403),
    .A(net408),
    .X(_0656_));
 sg13g2_nand2_1 _3604_ (.Y(_0657_),
    .A(_0638_),
    .B(_0656_));
 sg13g2_xnor2_1 _3605_ (.Y(_0658_),
    .A(_0638_),
    .B(_0656_));
 sg13g2_nor2_1 _3606_ (.A(_0654_),
    .B(_0658_),
    .Y(_0659_));
 sg13g2_and2_1 _3607_ (.A(net409),
    .B(net407),
    .X(_0660_));
 sg13g2_and3_2 _3608_ (.X(_0661_),
    .A(net409),
    .B(net408),
    .C(net407));
 sg13g2_a21oi_1 _3609_ (.A1(net409),
    .A2(net408),
    .Y(_0662_),
    .B1(net407));
 sg13g2_or2_1 _3610_ (.X(_0663_),
    .B(_0662_),
    .A(_0661_));
 sg13g2_inv_1 _3611_ (.Y(_0664_),
    .A(_0663_));
 sg13g2_xor2_1 _3612_ (.B(_0658_),
    .A(_0654_),
    .X(_0665_));
 sg13g2_a21oi_1 _3613_ (.A1(_0664_),
    .A2(_0665_),
    .Y(_0666_),
    .B1(_0659_));
 sg13g2_nand2_1 _3614_ (.Y(_0667_),
    .A(net409),
    .B(_0655_));
 sg13g2_inv_1 _3615_ (.Y(_0668_),
    .A(_0667_));
 sg13g2_xnor2_1 _3616_ (.Y(_0669_),
    .A(net409),
    .B(_0655_));
 sg13g2_inv_1 _3617_ (.Y(_0670_),
    .A(_0669_));
 sg13g2_xor2_1 _3618_ (.B(net403),
    .A(net405),
    .X(_0671_));
 sg13g2_nand2_1 _3619_ (.Y(_0672_),
    .A(_0640_),
    .B(_0671_));
 sg13g2_xnor2_1 _3620_ (.Y(_0673_),
    .A(_0640_),
    .B(_0671_));
 sg13g2_nor2_1 _3621_ (.A(_0657_),
    .B(_0673_),
    .Y(_0674_));
 sg13g2_xor2_1 _3622_ (.B(_0673_),
    .A(_0657_),
    .X(_0675_));
 sg13g2_xnor2_1 _3623_ (.Y(_0676_),
    .A(_0669_),
    .B(_0675_));
 sg13g2_nor2b_1 _3624_ (.A(_0666_),
    .B_N(_0676_),
    .Y(_0677_));
 sg13g2_xnor2_1 _3625_ (.Y(_0678_),
    .A(_0666_),
    .B(_0676_));
 sg13g2_a21o_2 _3626_ (.A2(_0678_),
    .A1(_0661_),
    .B1(_0677_),
    .X(_0679_));
 sg13g2_a21oi_1 _3627_ (.A1(_0670_),
    .A2(_0675_),
    .Y(_0680_),
    .B1(_0674_));
 sg13g2_nand2_1 _3628_ (.Y(_0681_),
    .A(net405),
    .B(_0655_));
 sg13g2_a21oi_1 _3629_ (.A1(net405),
    .A2(_0647_),
    .Y(_0682_),
    .B1(_0642_));
 sg13g2_a21o_1 _3630_ (.A2(_0655_),
    .A1(net405),
    .B1(_0682_),
    .X(_0683_));
 sg13g2_inv_1 _3631_ (.Y(_0684_),
    .A(_0683_));
 sg13g2_mux4_1 _3632_ (.S0(net547),
    .A0(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[10] ),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[10] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[10] ),
    .A3(net535),
    .S1(net545),
    .X(_0685_));
 sg13g2_nand2_1 _3633_ (.Y(_0686_),
    .A(net404),
    .B(_0685_));
 sg13g2_or2_1 _3634_ (.X(_0687_),
    .B(_0685_),
    .A(net404));
 sg13g2_xor2_1 _3635_ (.B(_0685_),
    .A(net405),
    .X(_0688_));
 sg13g2_nand2_1 _3636_ (.Y(_0689_),
    .A(net406),
    .B(_0688_));
 sg13g2_xnor2_1 _3637_ (.Y(_0690_),
    .A(net406),
    .B(_0688_));
 sg13g2_nor2_1 _3638_ (.A(_0672_),
    .B(_0690_),
    .Y(_0691_));
 sg13g2_xor2_1 _3639_ (.B(_0690_),
    .A(_0672_),
    .X(_0692_));
 sg13g2_xnor2_1 _3640_ (.Y(_0693_),
    .A(_0683_),
    .B(_0692_));
 sg13g2_nor2b_1 _3641_ (.A(_0680_),
    .B_N(_0693_),
    .Y(_0694_));
 sg13g2_xnor2_1 _3642_ (.Y(_0695_),
    .A(_0680_),
    .B(_0693_));
 sg13g2_xnor2_1 _3643_ (.Y(_0696_),
    .A(_0667_),
    .B(_0695_));
 sg13g2_nand2_1 _3644_ (.Y(_0697_),
    .A(_0679_),
    .B(_0696_));
 sg13g2_xnor2_1 _3645_ (.Y(_0698_),
    .A(_0679_),
    .B(_0696_));
 sg13g2_xor2_1 _3646_ (.B(net407),
    .A(net409),
    .X(_0699_));
 sg13g2_nand2_1 _3647_ (.Y(_0700_),
    .A(_0639_),
    .B(_0699_));
 sg13g2_xnor2_1 _3648_ (.Y(_0701_),
    .A(_0637_),
    .B(_0653_));
 sg13g2_nor2_1 _3649_ (.A(_0700_),
    .B(_0701_),
    .Y(_0702_));
 sg13g2_and2_1 _3650_ (.A(_0643_),
    .B(net406),
    .X(_0703_));
 sg13g2_nand2_1 _3651_ (.Y(_0704_),
    .A(net406),
    .B(_0660_));
 sg13g2_inv_1 _3652_ (.Y(_0705_),
    .A(_0704_));
 sg13g2_xnor2_1 _3653_ (.Y(_0706_),
    .A(net406),
    .B(_0660_));
 sg13g2_inv_1 _3654_ (.Y(_0707_),
    .A(_0706_));
 sg13g2_xor2_1 _3655_ (.B(_0701_),
    .A(_0700_),
    .X(_0708_));
 sg13g2_a21oi_1 _3656_ (.A1(_0707_),
    .A2(_0708_),
    .Y(_0709_),
    .B1(_0702_));
 sg13g2_xnor2_1 _3657_ (.Y(_0710_),
    .A(_0663_),
    .B(_0665_));
 sg13g2_nor2b_1 _3658_ (.A(_0709_),
    .B_N(_0710_),
    .Y(_0711_));
 sg13g2_xnor2_1 _3659_ (.Y(_0712_),
    .A(_0709_),
    .B(_0710_));
 sg13g2_a21o_1 _3660_ (.A2(_0712_),
    .A1(_0705_),
    .B1(_0711_),
    .X(_0713_));
 sg13g2_xor2_1 _3661_ (.B(_0678_),
    .A(_0661_),
    .X(_0714_));
 sg13g2_nor2_1 _3662_ (.A(_0713_),
    .B(_0714_),
    .Y(_0715_));
 sg13g2_xnor2_1 _3663_ (.Y(_0716_),
    .A(_0704_),
    .B(_0712_));
 sg13g2_xnor2_1 _3664_ (.Y(_0717_),
    .A(_0707_),
    .B(_0708_));
 sg13g2_nand2_1 _3665_ (.Y(_0718_),
    .A(_0640_),
    .B(net406));
 sg13g2_xnor2_1 _3666_ (.Y(_0719_),
    .A(_0639_),
    .B(_0699_));
 sg13g2_xnor2_1 _3667_ (.Y(_0720_),
    .A(_0640_),
    .B(_0703_));
 sg13g2_nor2_1 _3668_ (.A(_0719_),
    .B(_0720_),
    .Y(_0721_));
 sg13g2_a21oi_1 _3669_ (.A1(_0640_),
    .A2(_0703_),
    .Y(_0722_),
    .B1(_0721_));
 sg13g2_nor2_1 _3670_ (.A(_0717_),
    .B(_0722_),
    .Y(_0723_));
 sg13g2_and2_1 _3671_ (.A(_0638_),
    .B(_0640_),
    .X(_0724_));
 sg13g2_nor2b_1 _3672_ (.A(_0718_),
    .B_N(_0638_),
    .Y(_0725_));
 sg13g2_o21ai_1 _3673_ (.B1(_0644_),
    .Y(_0726_),
    .A1(_0637_),
    .A2(_0638_));
 sg13g2_nor2b_1 _3674_ (.A(_0640_),
    .B_N(_0726_),
    .Y(_0727_));
 sg13g2_o21ai_1 _3675_ (.B1(_0718_),
    .Y(_0728_),
    .A1(_0648_),
    .A2(_0724_));
 sg13g2_o21ai_1 _3676_ (.B1(_0637_),
    .Y(_0729_),
    .A1(_0638_),
    .A2(_0639_));
 sg13g2_o21ai_1 _3677_ (.B1(_0729_),
    .Y(_0730_),
    .A1(_0727_),
    .A2(_0728_));
 sg13g2_nor2_1 _3678_ (.A(_0645_),
    .B(_0703_),
    .Y(_0731_));
 sg13g2_xor2_1 _3679_ (.B(_0718_),
    .A(_0638_),
    .X(_0732_));
 sg13g2_nor3_1 _3680_ (.A(_0645_),
    .B(_0703_),
    .C(_0732_),
    .Y(_0733_));
 sg13g2_xnor2_1 _3681_ (.Y(_0734_),
    .A(_0731_),
    .B(_0732_));
 sg13g2_nand3_1 _3682_ (.B(_0730_),
    .C(_0731_),
    .A(_0725_),
    .Y(_0735_));
 sg13g2_xor2_1 _3683_ (.B(_0720_),
    .A(_0719_),
    .X(_0736_));
 sg13g2_nor2_1 _3684_ (.A(_0733_),
    .B(_0736_),
    .Y(_0737_));
 sg13g2_nand3_1 _3685_ (.B(_0639_),
    .C(_0724_),
    .A(_0637_),
    .Y(_0738_));
 sg13g2_nand2b_1 _3686_ (.Y(_0739_),
    .B(_0738_),
    .A_N(_0725_));
 sg13g2_a221oi_1 _3687_ (.B2(_0733_),
    .C1(_0739_),
    .B1(_0736_),
    .A1(_0730_),
    .Y(_0740_),
    .A2(_0734_));
 sg13g2_a221oi_1 _3688_ (.B2(_0737_),
    .C1(_0740_),
    .B1(_0735_),
    .A1(_0717_),
    .Y(_0741_),
    .A2(_0722_));
 sg13g2_or2_1 _3689_ (.X(_0742_),
    .B(_0741_),
    .A(_0723_));
 sg13g2_a22oi_1 _3690_ (.Y(_0743_),
    .B1(_0716_),
    .B2(_0742_),
    .A2(_0714_),
    .A1(_0713_));
 sg13g2_nor2_1 _3691_ (.A(_0715_),
    .B(_0743_),
    .Y(_0744_));
 sg13g2_nor3_1 _3692_ (.A(_0698_),
    .B(_0715_),
    .C(_0743_),
    .Y(_0745_));
 sg13g2_xor2_1 _3693_ (.B(_0744_),
    .A(_0698_),
    .X(_0746_));
 sg13g2_and2_1 _3694_ (.A(_0652_),
    .B(_0746_),
    .X(_0747_));
 sg13g2_a21oi_1 _3695_ (.A1(_0668_),
    .A2(_0695_),
    .Y(_0748_),
    .B1(_0694_));
 sg13g2_a21oi_1 _3696_ (.A1(_0684_),
    .A2(_0692_),
    .Y(_0749_),
    .B1(_0691_));
 sg13g2_nand3_1 _3697_ (.B(net403),
    .C(_0685_),
    .A(net404),
    .Y(_0750_));
 sg13g2_xor2_1 _3698_ (.B(_0686_),
    .A(net403),
    .X(_0751_));
 sg13g2_inv_1 _3699_ (.Y(_0752_),
    .A(_0751_));
 sg13g2_nand2_1 _3700_ (.Y(_0753_),
    .A(_0636_),
    .B(_0685_));
 sg13g2_xor2_1 _3701_ (.B(_0685_),
    .A(_0636_),
    .X(_0754_));
 sg13g2_inv_1 _3702_ (.Y(_0755_),
    .A(_0754_));
 sg13g2_xnor2_1 _3703_ (.Y(_0756_),
    .A(net407),
    .B(_0754_));
 sg13g2_nor2_1 _3704_ (.A(_0689_),
    .B(_0756_),
    .Y(_0757_));
 sg13g2_xor2_1 _3705_ (.B(_0756_),
    .A(_0689_),
    .X(_0758_));
 sg13g2_xnor2_1 _3706_ (.Y(_0759_),
    .A(_0751_),
    .B(_0758_));
 sg13g2_nand2b_1 _3707_ (.Y(_0760_),
    .B(_0759_),
    .A_N(_0749_));
 sg13g2_xnor2_1 _3708_ (.Y(_0761_),
    .A(_0749_),
    .B(_0759_));
 sg13g2_nand2b_1 _3709_ (.Y(_0762_),
    .B(_0761_),
    .A_N(_0681_));
 sg13g2_xnor2_1 _3710_ (.Y(_0763_),
    .A(_0681_),
    .B(_0761_));
 sg13g2_nor2b_1 _3711_ (.A(_0763_),
    .B_N(_0748_),
    .Y(_0764_));
 sg13g2_nand2b_1 _3712_ (.Y(_0765_),
    .B(_0763_),
    .A_N(_0748_));
 sg13g2_xor2_1 _3713_ (.B(_0763_),
    .A(_0748_),
    .X(_0766_));
 sg13g2_a21oi_1 _3714_ (.A1(_0679_),
    .A2(_0696_),
    .Y(_0767_),
    .B1(_0745_));
 sg13g2_xnor2_1 _3715_ (.Y(_0768_),
    .A(_0766_),
    .B(_0767_));
 sg13g2_nand2_1 _3716_ (.Y(_0769_),
    .A(_0747_),
    .B(_0768_));
 sg13g2_nor2_1 _3717_ (.A(_0698_),
    .B(_0766_),
    .Y(_0770_));
 sg13g2_a21oi_1 _3718_ (.A1(_0697_),
    .A2(_0765_),
    .Y(_0771_),
    .B1(_0764_));
 sg13g2_a21oi_2 _3719_ (.B1(_0771_),
    .Y(_0772_),
    .A2(_0770_),
    .A1(_0744_));
 sg13g2_nand2_1 _3720_ (.Y(_0773_),
    .A(_0760_),
    .B(_0762_));
 sg13g2_a21oi_1 _3721_ (.A1(_0752_),
    .A2(_0758_),
    .Y(_0774_),
    .B1(_0757_));
 sg13g2_nand3_1 _3722_ (.B(net404),
    .C(_0685_),
    .A(_0636_),
    .Y(_0775_));
 sg13g2_xor2_1 _3723_ (.B(_0753_),
    .A(net404),
    .X(_0776_));
 sg13g2_nand2_1 _3724_ (.Y(_0777_),
    .A(_0660_),
    .B(_0754_));
 sg13g2_a21o_1 _3725_ (.A2(_0754_),
    .A1(net407),
    .B1(net409),
    .X(_0778_));
 sg13g2_nand2_1 _3726_ (.Y(_0779_),
    .A(_0777_),
    .B(_0778_));
 sg13g2_xor2_1 _3727_ (.B(_0779_),
    .A(_0776_),
    .X(_0780_));
 sg13g2_nor2b_1 _3728_ (.A(_0774_),
    .B_N(_0780_),
    .Y(_0781_));
 sg13g2_xnor2_1 _3729_ (.Y(_0782_),
    .A(_0774_),
    .B(_0780_));
 sg13g2_nor2b_1 _3730_ (.A(_0750_),
    .B_N(_0782_),
    .Y(_0783_));
 sg13g2_xnor2_1 _3731_ (.Y(_0784_),
    .A(_0750_),
    .B(_0782_));
 sg13g2_nand2_1 _3732_ (.Y(_0785_),
    .A(_0773_),
    .B(_0784_));
 sg13g2_xnor2_1 _3733_ (.Y(_0786_),
    .A(_0773_),
    .B(_0784_));
 sg13g2_xnor2_1 _3734_ (.Y(_0787_),
    .A(_0772_),
    .B(_0786_));
 sg13g2_nand3_1 _3735_ (.B(_0768_),
    .C(_0787_),
    .A(_0747_),
    .Y(_0788_));
 sg13g2_o21ai_1 _3736_ (.B1(_0777_),
    .Y(_0789_),
    .A1(_0776_),
    .A2(_0779_));
 sg13g2_nand2_1 _3737_ (.Y(_0790_),
    .A(net408),
    .B(_0754_));
 sg13g2_xnor2_1 _3738_ (.Y(_0791_),
    .A(net408),
    .B(_0754_));
 sg13g2_nand2b_1 _3739_ (.Y(_0792_),
    .B(_0789_),
    .A_N(_0791_));
 sg13g2_xor2_1 _3740_ (.B(_0791_),
    .A(_0789_),
    .X(_0793_));
 sg13g2_xor2_1 _3741_ (.B(_0793_),
    .A(_0775_),
    .X(_0794_));
 sg13g2_nor3_1 _3742_ (.A(_0781_),
    .B(_0783_),
    .C(_0794_),
    .Y(_0795_));
 sg13g2_o21ai_1 _3743_ (.B1(_0794_),
    .Y(_0796_),
    .A1(_0781_),
    .A2(_0783_));
 sg13g2_nor2b_1 _3744_ (.A(_0795_),
    .B_N(_0796_),
    .Y(_0797_));
 sg13g2_o21ai_1 _3745_ (.B1(_0785_),
    .Y(_0798_),
    .A1(_0772_),
    .A2(_0786_));
 sg13g2_xor2_1 _3746_ (.B(_0798_),
    .A(_0797_),
    .X(_0799_));
 sg13g2_o21ai_1 _3747_ (.B1(_0792_),
    .Y(_0800_),
    .A1(_0775_),
    .A2(_0793_));
 sg13g2_nand2_1 _3748_ (.Y(_0801_),
    .A(_0753_),
    .B(_0790_));
 sg13g2_nand2_1 _3749_ (.Y(_0802_),
    .A(net403),
    .B(_0801_));
 sg13g2_inv_1 _3750_ (.Y(_0803_),
    .A(_0802_));
 sg13g2_xor2_1 _3751_ (.B(_0801_),
    .A(net403),
    .X(_0804_));
 sg13g2_and2_1 _3752_ (.A(_0800_),
    .B(_0804_),
    .X(_0805_));
 sg13g2_xnor2_1 _3753_ (.Y(_0806_),
    .A(_0800_),
    .B(_0804_));
 sg13g2_inv_1 _3754_ (.Y(_0807_),
    .A(_0806_));
 sg13g2_nand2b_1 _3755_ (.Y(_0808_),
    .B(_0797_),
    .A_N(_0786_));
 sg13g2_a21o_1 _3756_ (.A2(_0796_),
    .A1(_0785_),
    .B1(_0795_),
    .X(_0809_));
 sg13g2_o21ai_1 _3757_ (.B1(_0809_),
    .Y(_0810_),
    .A1(_0772_),
    .A2(_0808_));
 sg13g2_xnor2_1 _3758_ (.Y(_0811_),
    .A(_0806_),
    .B(_0810_));
 sg13g2_o21ai_1 _3759_ (.B1(_0811_),
    .Y(_0812_),
    .A1(_0788_),
    .A2(_0799_));
 sg13g2_xor2_1 _3760_ (.B(net404),
    .A(_0636_),
    .X(_0813_));
 sg13g2_xnor2_1 _3761_ (.Y(_0814_),
    .A(_0802_),
    .B(_0813_));
 sg13g2_a21oi_1 _3762_ (.A1(_0807_),
    .A2(_0810_),
    .Y(_0815_),
    .B1(_0805_));
 sg13g2_xor2_1 _3763_ (.B(_0815_),
    .A(_0814_),
    .X(_0816_));
 sg13g2_or2_1 _3764_ (.X(_0817_),
    .B(_0816_),
    .A(_0812_));
 sg13g2_a21oi_1 _3765_ (.A1(_0812_),
    .A2(_0816_),
    .Y(_0818_),
    .B1(_0539_));
 sg13g2_a22oi_1 _3766_ (.Y(_0004_),
    .B1(_0817_),
    .B2(_0818_),
    .A2(_0551_),
    .A1(_0539_));
 sg13g2_nor2b_1 _3767_ (.A(net553),
    .B_N(net835),
    .Y(_0005_));
 sg13g2_nor2b_1 _3768_ (.A(net553),
    .B_N(net813),
    .Y(_0006_));
 sg13g2_nor2_1 _3769_ (.A(net419),
    .B(net792),
    .Y(_0007_));
 sg13g2_o21ai_1 _3770_ (.B1(net441),
    .Y(_0819_),
    .A1(net792),
    .A2(net831));
 sg13g2_a21oi_1 _3771_ (.A1(net792),
    .A2(net831),
    .Y(_0008_),
    .B1(_0819_));
 sg13g2_nand2_1 _3772_ (.Y(_0820_),
    .A(_0539_),
    .B(net895));
 sg13g2_nor4_1 _3773_ (.A(_0542_),
    .B(net936),
    .C(net950),
    .D(net874),
    .Y(_0821_));
 sg13g2_or3_1 _3774_ (.A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[10] ),
    .B(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[9] ),
    .C(_0540_),
    .X(_0822_));
 sg13g2_nor4_1 _3775_ (.A(net1019),
    .B(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[5] ),
    .C(net1023),
    .D(_0822_),
    .Y(_0823_));
 sg13g2_nand4_1 _3776_ (.B(net941),
    .C(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[5] ),
    .A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[7] ),
    .Y(_0824_),
    .D(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[4] ));
 sg13g2_nor4_1 _3777_ (.A(net978),
    .B(net920),
    .C(net1024),
    .D(_0824_),
    .Y(_0825_));
 sg13g2_a21oi_1 _3778_ (.A1(_0821_),
    .A2(_0823_),
    .Y(_0826_),
    .B1(_0825_));
 sg13g2_a21oi_1 _3779_ (.A1(_0540_),
    .A2(_0541_),
    .Y(_0827_),
    .B1(_0627_));
 sg13g2_nor4_1 _3780_ (.A(net863),
    .B(net1001),
    .C(net983),
    .D(_0827_),
    .Y(_0828_));
 sg13g2_nand3b_1 _3781_ (.B(_0828_),
    .C(net554),
    .Y(_0829_),
    .A_N(_0630_));
 sg13g2_o21ai_1 _3782_ (.B1(net896),
    .Y(_0009_),
    .A1(_0826_),
    .A2(_0829_));
 sg13g2_nor2b_1 _3783_ (.A(net554),
    .B_N(net1065),
    .Y(_0830_));
 sg13g2_nand2b_1 _3784_ (.Y(_0831_),
    .B(net944),
    .A_N(net1003));
 sg13g2_a22oi_1 _3785_ (.Y(_0832_),
    .B1(_0549_),
    .B2(net978),
    .A2(_0548_),
    .A1(net920));
 sg13g2_nand2b_1 _3786_ (.Y(_0833_),
    .B(net929),
    .A_N(net1056));
 sg13g2_xor2_1 _3787_ (.B(net869),
    .A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[7] ),
    .X(_0834_));
 sg13g2_xor2_1 _3788_ (.B(net906),
    .A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[1] ),
    .X(_0835_));
 sg13g2_a221oi_1 _3789_ (.B2(net914),
    .C1(_0835_),
    .B1(_0552_),
    .A1(_0535_),
    .Y(_0836_),
    .A2(net909));
 sg13g2_a221oi_1 _3790_ (.B2(_0534_),
    .C1(_0834_),
    .B1(net889),
    .A1(net1003),
    .Y(_0837_),
    .A2(_0550_));
 sg13g2_xnor2_1 _3791_ (.Y(_0838_),
    .A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[9] ),
    .B(net835));
 sg13g2_xor2_1 _3792_ (.B(net882),
    .A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[0] ),
    .X(_0839_));
 sg13g2_xor2_1 _3793_ (.B(net866),
    .A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[6] ),
    .X(_0840_));
 sg13g2_nor4_1 _3794_ (.A(net863),
    .B(net813),
    .C(_0839_),
    .D(_0840_),
    .Y(_0841_));
 sg13g2_nand4_1 _3795_ (.B(_0837_),
    .C(_0838_),
    .A(_0836_),
    .Y(_0842_),
    .D(_0841_));
 sg13g2_a22oi_1 _3796_ (.Y(_0843_),
    .B1(_0551_),
    .B2(net1056),
    .A2(net892),
    .A1(_0536_));
 sg13g2_nand4_1 _3797_ (.B(_0832_),
    .C(_0833_),
    .A(_0831_),
    .Y(_0844_),
    .D(_0843_));
 sg13g2_nor3_1 _3798_ (.A(_0829_),
    .B(_0842_),
    .C(_0844_),
    .Y(_0845_));
 sg13g2_a21o_1 _3799_ (.A2(_0845_),
    .A1(_0826_),
    .B1(net1066),
    .X(_0010_));
 sg13g2_o21ai_1 _3800_ (.B1(net451),
    .Y(_0846_),
    .A1(_0651_),
    .A2(_0685_));
 sg13g2_nor2_1 _3801_ (.A(_0636_),
    .B(_0846_),
    .Y(_0011_));
 sg13g2_xnor2_1 _3802_ (.Y(_0847_),
    .A(_0652_),
    .B(_0746_));
 sg13g2_nor2_1 _3803_ (.A(net553),
    .B(net882),
    .Y(_0848_));
 sg13g2_a21oi_1 _3804_ (.A1(net553),
    .A2(_0847_),
    .Y(_0012_),
    .B1(net883));
 sg13g2_nor2_1 _3805_ (.A(net552),
    .B(net906),
    .Y(_0849_));
 sg13g2_xnor2_1 _3806_ (.Y(_0850_),
    .A(_0747_),
    .B(_0768_));
 sg13g2_a21oi_1 _3807_ (.A1(net552),
    .A2(_0850_),
    .Y(_0013_),
    .B1(net907));
 sg13g2_xor2_1 _3808_ (.B(_0787_),
    .A(_0769_),
    .X(_0851_));
 sg13g2_nor2_1 _3809_ (.A(net553),
    .B(net892),
    .Y(_0852_));
 sg13g2_a21oi_1 _3810_ (.A1(net552),
    .A2(_0851_),
    .Y(_0014_),
    .B1(net893));
 sg13g2_nor2_1 _3811_ (.A(net552),
    .B(net909),
    .Y(_0853_));
 sg13g2_xnor2_1 _3812_ (.Y(_0854_),
    .A(_0788_),
    .B(_0799_));
 sg13g2_a21oi_1 _3813_ (.A1(net552),
    .A2(_0854_),
    .Y(_0015_),
    .B1(net910));
 sg13g2_or3_1 _3814_ (.A(_0788_),
    .B(_0799_),
    .C(_0811_),
    .X(_0855_));
 sg13g2_and2_1 _3815_ (.A(net552),
    .B(_0812_),
    .X(_0856_));
 sg13g2_a22oi_1 _3816_ (.Y(_0016_),
    .B1(_0855_),
    .B2(_0856_),
    .A2(_0550_),
    .A1(_0539_));
 sg13g2_nor2_1 _3817_ (.A(net553),
    .B(net866),
    .Y(_0857_));
 sg13g2_o21ai_1 _3818_ (.B1(_0813_),
    .Y(_0858_),
    .A1(_0803_),
    .A2(_0805_));
 sg13g2_nand2_1 _3819_ (.Y(_0859_),
    .A(_0807_),
    .B(_0814_));
 sg13g2_o21ai_1 _3820_ (.B1(_0858_),
    .Y(_0860_),
    .A1(_0809_),
    .A2(_0859_));
 sg13g2_nor3_1 _3821_ (.A(_0772_),
    .B(_0808_),
    .C(_0859_),
    .Y(_0861_));
 sg13g2_or2_1 _3822_ (.X(_0862_),
    .B(_0861_),
    .A(_0860_));
 sg13g2_o21ai_1 _3823_ (.B1(_0686_),
    .Y(_0863_),
    .A1(net404),
    .A2(_0755_));
 sg13g2_xnor2_1 _3824_ (.Y(_0864_),
    .A(_0862_),
    .B(_0863_));
 sg13g2_nor3_1 _3825_ (.A(_0812_),
    .B(_0816_),
    .C(_0864_),
    .Y(_0865_));
 sg13g2_o21ai_1 _3826_ (.B1(_0864_),
    .Y(_0866_),
    .A1(_0812_),
    .A2(_0816_));
 sg13g2_nand3b_1 _3827_ (.B(_0866_),
    .C(net552),
    .Y(_0867_),
    .A_N(_0865_));
 sg13g2_nor2b_1 _3828_ (.A(net867),
    .B_N(_0867_),
    .Y(_0017_));
 sg13g2_nor2_1 _3829_ (.A(net553),
    .B(net869),
    .Y(_0868_));
 sg13g2_a22oi_1 _3830_ (.Y(_0869_),
    .B1(_0862_),
    .B2(_0863_),
    .A2(_0687_),
    .A1(_0636_));
 sg13g2_nor2b_1 _3831_ (.A(_0869_),
    .B_N(_0865_),
    .Y(_0870_));
 sg13g2_xnor2_1 _3832_ (.Y(_0871_),
    .A(_0865_),
    .B(_0869_));
 sg13g2_a21oi_1 _3833_ (.A1(net553),
    .A2(_0871_),
    .Y(_0018_),
    .B1(net870));
 sg13g2_nand2_1 _3834_ (.Y(_0872_),
    .A(_0539_),
    .B(net889));
 sg13g2_nand2_1 _3835_ (.Y(_0873_),
    .A(net552),
    .B(_0636_));
 sg13g2_o21ai_1 _3836_ (.B1(net890),
    .Y(_0019_),
    .A1(_0870_),
    .A2(_0873_));
 sg13g2_o21ai_1 _3837_ (.B1(net441),
    .Y(_0874_),
    .A1(net554),
    .A2(net857));
 sg13g2_a21oi_1 _3838_ (.A1(net554),
    .A2(net857),
    .Y(_0020_),
    .B1(_0874_));
 sg13g2_a21oi_1 _3839_ (.A1(net554),
    .A2(net857),
    .Y(_0875_),
    .B1(net874));
 sg13g2_and3_1 _3840_ (.X(_0876_),
    .A(net554),
    .B(net874),
    .C(net857));
 sg13g2_nor3_1 _3841_ (.A(net419),
    .B(net875),
    .C(_0876_),
    .Y(_0021_));
 sg13g2_nor2_1 _3842_ (.A(net950),
    .B(_0876_),
    .Y(_0877_));
 sg13g2_and2_1 _3843_ (.A(net950),
    .B(_0876_),
    .X(_0878_));
 sg13g2_nor3_1 _3844_ (.A(net419),
    .B(net951),
    .C(_0878_),
    .Y(_0022_));
 sg13g2_nor2_1 _3845_ (.A(net936),
    .B(_0878_),
    .Y(_0879_));
 sg13g2_and2_1 _3846_ (.A(net936),
    .B(_0878_),
    .X(_0880_));
 sg13g2_nor3_1 _3847_ (.A(net419),
    .B(net937),
    .C(_0880_),
    .Y(_0023_));
 sg13g2_and2_1 _3848_ (.A(net1023),
    .B(_0880_),
    .X(_0881_));
 sg13g2_o21ai_1 _3849_ (.B1(net441),
    .Y(_0882_),
    .A1(net1023),
    .A2(_0880_));
 sg13g2_nor2_1 _3850_ (.A(_0881_),
    .B(_0882_),
    .Y(_0024_));
 sg13g2_nor3_1 _3851_ (.A(net1019),
    .B(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[6] ),
    .C(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[5] ),
    .Y(_0883_));
 sg13g2_and3_2 _3852_ (.X(_0884_),
    .A(_0827_),
    .B(_0881_),
    .C(_0883_));
 sg13g2_nor2_2 _3853_ (.A(net419),
    .B(_0884_),
    .Y(_0885_));
 sg13g2_and2_1 _3854_ (.A(net1040),
    .B(_0881_),
    .X(_0886_));
 sg13g2_o21ai_1 _3855_ (.B1(_0885_),
    .Y(_0887_),
    .A1(net1040),
    .A2(_0881_));
 sg13g2_nor2_1 _3856_ (.A(_0886_),
    .B(_0887_),
    .Y(_0025_));
 sg13g2_and2_1 _3857_ (.A(net1030),
    .B(_0886_),
    .X(_0888_));
 sg13g2_o21ai_1 _3858_ (.B1(net441),
    .Y(_0889_),
    .A1(net1030),
    .A2(_0886_));
 sg13g2_nor2_1 _3859_ (.A(_0888_),
    .B(net1031),
    .Y(_0026_));
 sg13g2_and2_1 _3860_ (.A(net1019),
    .B(_0888_),
    .X(_0890_));
 sg13g2_o21ai_1 _3861_ (.B1(net441),
    .Y(_0891_),
    .A1(net1019),
    .A2(_0888_));
 sg13g2_nor2_1 _3862_ (.A(_0890_),
    .B(net1020),
    .Y(_0027_));
 sg13g2_o21ai_1 _3863_ (.B1(_0885_),
    .Y(_0892_),
    .A1(net842),
    .A2(_0890_));
 sg13g2_a21oi_1 _3864_ (.A1(net842),
    .A2(_0890_),
    .Y(_0028_),
    .B1(_0892_));
 sg13g2_a21oi_1 _3865_ (.A1(net842),
    .A2(_0890_),
    .Y(_0893_),
    .B1(net887));
 sg13g2_nand3_1 _3866_ (.B(net842),
    .C(_0890_),
    .A(net887),
    .Y(_0894_));
 sg13g2_nand2_1 _3867_ (.Y(_0895_),
    .A(_0885_),
    .B(_0894_));
 sg13g2_nor2_1 _3868_ (.A(net888),
    .B(_0895_),
    .Y(_0029_));
 sg13g2_o21ai_1 _3869_ (.B1(net441),
    .Y(_0896_),
    .A1(_0538_),
    .A2(_0894_));
 sg13g2_a21oi_1 _3870_ (.A1(_0538_),
    .A2(_0894_),
    .Y(_0030_),
    .B1(_0896_));
 sg13g2_nor3_1 _3871_ (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[6] ),
    .B(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[5] ),
    .C(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[0] ),
    .Y(_0897_));
 sg13g2_nor3_1 _3872_ (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[10] ),
    .B(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[8] ),
    .C(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[7] ),
    .Y(_0898_));
 sg13g2_nor3_1 _3873_ (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[4] ),
    .B(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[1] ),
    .C(_0632_),
    .Y(_0899_));
 sg13g2_nand4_1 _3874_ (.B(_0897_),
    .C(_0898_),
    .A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[9] ),
    .Y(_0900_),
    .D(_0899_));
 sg13g2_and2_1 _3875_ (.A(_0884_),
    .B(_0900_),
    .X(_0901_));
 sg13g2_nand2_1 _3876_ (.Y(_0902_),
    .A(net1093),
    .B(_0884_));
 sg13g2_o21ai_1 _3877_ (.B1(_0902_),
    .Y(_0903_),
    .A1(net1093),
    .A2(_0901_));
 sg13g2_nor2_1 _3878_ (.A(net419),
    .B(net1094),
    .Y(_0031_));
 sg13g2_nand2_1 _3879_ (.Y(_0904_),
    .A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[1] ),
    .B(net1577));
 sg13g2_o21ai_1 _3880_ (.B1(net443),
    .Y(_0905_),
    .A1(_0537_),
    .A2(_0902_));
 sg13g2_a21oi_1 _3881_ (.A1(_0537_),
    .A2(_0902_),
    .Y(_0032_),
    .B1(_0905_));
 sg13g2_nand2_1 _3882_ (.Y(_0906_),
    .A(net920),
    .B(_0885_));
 sg13g2_nand3_1 _3883_ (.B(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[1] ),
    .C(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[0] ),
    .A(net920),
    .Y(_0907_));
 sg13g2_xnor2_1 _3884_ (.Y(_0908_),
    .A(_0536_),
    .B(_0904_));
 sg13g2_nand2_1 _3885_ (.Y(_0909_),
    .A(net443),
    .B(_0901_));
 sg13g2_o21ai_1 _3886_ (.B1(_0906_),
    .Y(_0033_),
    .A1(_0908_),
    .A2(_0909_));
 sg13g2_and2_1 _3887_ (.A(_0535_),
    .B(_0907_),
    .X(_0910_));
 sg13g2_nor2_2 _3888_ (.A(_0632_),
    .B(_0904_),
    .Y(_0911_));
 sg13g2_nor3_1 _3889_ (.A(_0909_),
    .B(_0910_),
    .C(_0911_),
    .Y(_0912_));
 sg13g2_a21o_1 _3890_ (.A2(_0885_),
    .A1(net978),
    .B1(_0912_),
    .X(_0034_));
 sg13g2_a21oi_1 _3891_ (.A1(_0884_),
    .A2(_0911_),
    .Y(_0913_),
    .B1(net1003));
 sg13g2_nand3_1 _3892_ (.B(_0884_),
    .C(_0911_),
    .A(net1003),
    .Y(_0914_));
 sg13g2_inv_1 _3893_ (.Y(_0915_),
    .A(_0914_));
 sg13g2_nor3_1 _3894_ (.A(net420),
    .B(net1004),
    .C(_0915_),
    .Y(_0035_));
 sg13g2_xor2_1 _3895_ (.B(_0914_),
    .A(net1056),
    .X(_0916_));
 sg13g2_nor2_1 _3896_ (.A(net420),
    .B(_0916_),
    .Y(_0036_));
 sg13g2_a21oi_1 _3897_ (.A1(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[5] ),
    .A2(_0915_),
    .Y(_0917_),
    .B1(net941));
 sg13g2_and3_2 _3898_ (.X(_0918_),
    .A(net941),
    .B(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[5] ),
    .C(_0915_));
 sg13g2_nor3_1 _3899_ (.A(net420),
    .B(net942),
    .C(_0918_),
    .Y(_0037_));
 sg13g2_o21ai_1 _3900_ (.B1(net443),
    .Y(_0919_),
    .A1(net901),
    .A2(_0918_));
 sg13g2_a21oi_1 _3901_ (.A1(net901),
    .A2(_0918_),
    .Y(_0038_),
    .B1(_0919_));
 sg13g2_a21oi_1 _3902_ (.A1(net901),
    .A2(_0918_),
    .Y(_0920_),
    .B1(net914));
 sg13g2_nand3_1 _3903_ (.B(_0630_),
    .C(_0911_),
    .A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[4] ),
    .Y(_0921_));
 sg13g2_and2_1 _3904_ (.A(_0630_),
    .B(_0915_),
    .X(_0922_));
 sg13g2_nor3_1 _3905_ (.A(net420),
    .B(net915),
    .C(_0922_),
    .Y(_0039_));
 sg13g2_nand2_1 _3906_ (.Y(_0923_),
    .A(net1001),
    .B(_0885_));
 sg13g2_xor2_1 _3907_ (.B(_0921_),
    .A(net1001),
    .X(_0924_));
 sg13g2_o21ai_1 _3908_ (.B1(_0923_),
    .Y(_0040_),
    .A1(_0909_),
    .A2(_0924_));
 sg13g2_and2_1 _3909_ (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[9] ),
    .B(_0922_),
    .X(_0925_));
 sg13g2_o21ai_1 _3910_ (.B1(net443),
    .Y(_0926_),
    .A1(net863),
    .A2(_0925_));
 sg13g2_a21oi_1 _3911_ (.A1(net863),
    .A2(_0925_),
    .Y(_0041_),
    .B1(_0926_));
 sg13g2_and3_1 _3912_ (.X(_0042_),
    .A(net441),
    .B(net792),
    .C(net831));
 sg13g2_and2_1 _3913_ (.A(net469),
    .B(net800),
    .X(_0043_));
 sg13g2_and2_1 _3914_ (.A(net464),
    .B(net774),
    .X(_0044_));
 sg13g2_and2_1 _3915_ (.A(net463),
    .B(net790),
    .X(_0045_));
 sg13g2_and2_1 _3916_ (.A(net463),
    .B(net820),
    .X(_0046_));
 sg13g2_and2_1 _3917_ (.A(net463),
    .B(net805),
    .X(_0047_));
 sg13g2_and2_1 _3918_ (.A(net463),
    .B(net808),
    .X(_0048_));
 sg13g2_and2_1 _3919_ (.A(net450),
    .B(net781),
    .X(_0049_));
 sg13g2_and2_1 _3920_ (.A(net450),
    .B(net776),
    .X(_0050_));
 sg13g2_and2_1 _3921_ (.A(net465),
    .B(net807),
    .X(_0051_));
 sg13g2_and2_1 _3922_ (.A(net463),
    .B(net788),
    .X(_0052_));
 sg13g2_and2_1 _3923_ (.A(net463),
    .B(net795),
    .X(_0053_));
 sg13g2_and2_1 _3924_ (.A(net464),
    .B(net825),
    .X(_0054_));
 sg13g2_and2_1 _3925_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[1] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[0] ),
    .X(_0927_));
 sg13g2_nor3_1 _3926_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[3] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[2] ),
    .C(_0927_),
    .Y(_0928_));
 sg13g2_nor2b_1 _3927_ (.A(_0928_),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[4] ),
    .Y(_0929_));
 sg13g2_o21ai_1 _3928_ (.B1(net952),
    .Y(_0930_),
    .A1(net961),
    .A2(_0929_));
 sg13g2_nand4_1 _3929_ (.B(net982),
    .C(net1012),
    .A(_0532_),
    .Y(_0931_),
    .D(net918));
 sg13g2_a21oi_1 _3930_ (.A1(_0533_),
    .A2(_0930_),
    .Y(_0932_),
    .B1(_0931_));
 sg13g2_or2_1 _3931_ (.X(_0933_),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[0] ),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[1] ));
 sg13g2_nand3_1 _3932_ (.B(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[2] ),
    .C(_0933_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[3] ),
    .Y(_0934_));
 sg13g2_nand2b_1 _3933_ (.Y(_0935_),
    .B(_0934_),
    .A_N(net948));
 sg13g2_a21oi_1 _3934_ (.A1(net961),
    .A2(_0935_),
    .Y(_0936_),
    .B1(net952));
 sg13g2_nand2b_1 _3935_ (.Y(_0937_),
    .B(net885),
    .A_N(net548));
 sg13g2_nor4_1 _3936_ (.A(_0532_),
    .B(net982),
    .C(net1012),
    .D(net918),
    .Y(_0938_));
 sg13g2_nand2b_1 _3937_ (.Y(_0939_),
    .B(net918),
    .A_N(net548));
 sg13g2_or2_1 _3938_ (.X(_0940_),
    .B(_0938_),
    .A(net551));
 sg13g2_o21ai_1 _3939_ (.B1(_0940_),
    .Y(_0941_),
    .A1(_0936_),
    .A2(_0937_));
 sg13g2_o21ai_1 _3940_ (.B1(net450),
    .Y(_0055_),
    .A1(_0932_),
    .A2(_0941_));
 sg13g2_nor3_1 _3941_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt_sum[5] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[1] ),
    .C(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[2] ),
    .Y(_0942_));
 sg13g2_or4_1 _3942_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt_sum[5] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[1] ),
    .C(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[2] ),
    .D(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[3] ),
    .X(_0943_));
 sg13g2_nor3_1 _3943_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[4] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[5] ),
    .C(_0943_),
    .Y(_0944_));
 sg13g2_nor2b_1 _3944_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[6] ),
    .B_N(_0944_),
    .Y(_0945_));
 sg13g2_nand2b_2 _3945_ (.Y(_0946_),
    .B(_0945_),
    .A_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[7] ));
 sg13g2_nor3_1 _3946_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[8] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[9] ),
    .C(_0946_),
    .Y(_0947_));
 sg13g2_nor2b_1 _3947_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[10] ),
    .B_N(_0947_),
    .Y(_0948_));
 sg13g2_xor2_1 _3948_ (.B(_0946_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[8] ),
    .X(_0949_));
 sg13g2_xnor2_1 _3949_ (.Y(_0950_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[13] ),
    .B(_0949_));
 sg13g2_xor2_1 _3950_ (.B(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[17] ),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[12] ),
    .X(_0951_));
 sg13g2_o21ai_1 _3951_ (.B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[9] ),
    .Y(_0952_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[8] ),
    .A2(_0946_));
 sg13g2_nor2b_1 _3952_ (.A(_0947_),
    .B_N(_0952_),
    .Y(_0953_));
 sg13g2_xnor2_1 _3953_ (.Y(_0954_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[14] ),
    .B(_0953_));
 sg13g2_xnor2_1 _3954_ (.Y(_0955_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[4] ),
    .B(_0943_));
 sg13g2_o21ai_1 _3955_ (.B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[2] ),
    .Y(_0956_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt_sum[5] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[1] ));
 sg13g2_nor2b_1 _3956_ (.A(_0942_),
    .B_N(_0956_),
    .Y(_0957_));
 sg13g2_nor2_1 _3957_ (.A(net763),
    .B(net1007),
    .Y(_0958_));
 sg13g2_xnor2_1 _3958_ (.Y(_0959_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[5] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt_sum[5] ));
 sg13g2_nand2_1 _3959_ (.Y(_0960_),
    .A(_0958_),
    .B(_0959_));
 sg13g2_nor4_1 _3960_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[3] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[2] ),
    .C(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[4] ),
    .D(_0960_),
    .Y(_0961_));
 sg13g2_o21ai_1 _3961_ (.B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[5] ),
    .Y(_0962_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[4] ),
    .A2(_0943_));
 sg13g2_nor2b_1 _3962_ (.A(_0944_),
    .B_N(_0962_),
    .Y(_0963_));
 sg13g2_xnor2_1 _3963_ (.Y(_0964_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[3] ),
    .B(_0942_));
 sg13g2_xor2_1 _3964_ (.B(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[1] ),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt_sum[5] ),
    .X(_0965_));
 sg13g2_xnor2_1 _3965_ (.Y(_0966_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[6] ),
    .B(_0965_));
 sg13g2_xnor2_1 _3966_ (.Y(_0967_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[7] ),
    .B(_0945_));
 sg13g2_xor2_1 _3967_ (.B(_0944_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[6] ),
    .X(_0968_));
 sg13g2_xnor2_1 _3968_ (.Y(_0969_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[11] ),
    .B(_0968_));
 sg13g2_xnor2_1 _3969_ (.Y(_0970_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[7] ),
    .B(_0957_));
 sg13g2_xnor2_1 _3970_ (.Y(_0971_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[8] ),
    .B(_0964_));
 sg13g2_nand4_1 _3971_ (.B(_0966_),
    .C(_0970_),
    .A(_0961_),
    .Y(_0972_),
    .D(_0971_));
 sg13g2_xnor2_1 _3972_ (.Y(_0973_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[9] ),
    .B(_0955_));
 sg13g2_xor2_1 _3973_ (.B(_0963_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[10] ),
    .X(_0974_));
 sg13g2_nor4_1 _3974_ (.A(_0969_),
    .B(_0972_),
    .C(_0973_),
    .D(_0974_),
    .Y(_0975_));
 sg13g2_xnor2_1 _3975_ (.Y(_0976_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[12] ),
    .B(_0967_));
 sg13g2_nand4_1 _3976_ (.B(_0954_),
    .C(_0975_),
    .A(_0950_),
    .Y(_0977_),
    .D(_0976_));
 sg13g2_nor2b_1 _3977_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[11] ),
    .B_N(_0948_),
    .Y(_0978_));
 sg13g2_xnor2_1 _3978_ (.Y(_0979_),
    .A(_0951_),
    .B(_0978_));
 sg13g2_xnor2_1 _3979_ (.Y(_0980_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[10] ),
    .B(_0947_));
 sg13g2_xnor2_1 _3980_ (.Y(_0981_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[15] ),
    .B(_0980_));
 sg13g2_nand2_1 _3981_ (.Y(_0982_),
    .A(_0979_),
    .B(_0981_));
 sg13g2_xnor2_1 _3982_ (.Y(_0983_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[11] ),
    .B(_0948_));
 sg13g2_nor2b_2 _3983_ (.A(_0983_),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[16] ),
    .Y(_0984_));
 sg13g2_nor2b_2 _3984_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[16] ),
    .B_N(_0983_),
    .Y(_0985_));
 sg13g2_nor4_2 _3985_ (.A(_0977_),
    .B(_0982_),
    .C(_0984_),
    .Y(_0986_),
    .D(_0985_));
 sg13g2_nor4_2 _3986_ (.A(_0977_),
    .B(_0982_),
    .C(_0984_),
    .Y(_0987_),
    .D(_0985_));
 sg13g2_nor2_1 _3987_ (.A(net423),
    .B(_0987_),
    .Y(_0988_));
 sg13g2_nand2b_1 _3988_ (.Y(_0989_),
    .B(net449),
    .A_N(_0987_));
 sg13g2_nand2_1 _3989_ (.Y(_0990_),
    .A(net940),
    .B(net377));
 sg13g2_nand2_1 _3990_ (.Y(_0991_),
    .A(net448),
    .B(_0986_));
 sg13g2_inv_2 _3991_ (.Y(_0992_),
    .A(net372));
 sg13g2_o21ai_1 _3992_ (.B1(_0990_),
    .Y(_0056_),
    .A1(net940),
    .A2(net372));
 sg13g2_nand2_1 _3993_ (.Y(_0993_),
    .A(net924),
    .B(net376));
 sg13g2_nand2_1 _3994_ (.Y(_0994_),
    .A(net924),
    .B(net549));
 sg13g2_xor2_1 _3995_ (.B(net550),
    .A(net924),
    .X(_0995_));
 sg13g2_and2_1 _3996_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[0] ),
    .B(_0995_),
    .X(_0996_));
 sg13g2_nand2_1 _3997_ (.Y(_0997_),
    .A(net940),
    .B(_0995_));
 sg13g2_o21ai_1 _3998_ (.B1(_0992_),
    .Y(_0998_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[0] ),
    .A2(_0995_));
 sg13g2_o21ai_1 _3999_ (.B1(_0993_),
    .Y(_0057_),
    .A1(_0996_),
    .A2(_0998_));
 sg13g2_nand2_1 _4000_ (.Y(_0999_),
    .A(net980),
    .B(net376));
 sg13g2_xnor2_1 _4001_ (.Y(_1000_),
    .A(net980),
    .B(net550));
 sg13g2_a21oi_1 _4002_ (.A1(_0994_),
    .A2(_0997_),
    .Y(_1001_),
    .B1(_1000_));
 sg13g2_nand3_1 _4003_ (.B(_0997_),
    .C(_1000_),
    .A(_0994_),
    .Y(_1002_));
 sg13g2_nand2b_1 _4004_ (.Y(_1003_),
    .B(_1002_),
    .A_N(_1001_));
 sg13g2_o21ai_1 _4005_ (.B1(_0999_),
    .Y(_0058_),
    .A1(net372),
    .A2(_1003_));
 sg13g2_nand2_1 _4006_ (.Y(_1004_),
    .A(net954),
    .B(net376));
 sg13g2_a21oi_1 _4007_ (.A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[2] ),
    .A2(net549),
    .Y(_1005_),
    .B1(_1001_));
 sg13g2_nor2_1 _4008_ (.A(net954),
    .B(net550),
    .Y(_1006_));
 sg13g2_nand2_1 _4009_ (.Y(_1007_),
    .A(net954),
    .B(net549));
 sg13g2_nand2b_1 _4010_ (.Y(_1008_),
    .B(_1007_),
    .A_N(_1006_));
 sg13g2_xnor2_1 _4011_ (.Y(_1009_),
    .A(_1005_),
    .B(_1008_));
 sg13g2_o21ai_1 _4012_ (.B1(_1004_),
    .Y(_0059_),
    .A1(net372),
    .A2(_1009_));
 sg13g2_nand2_1 _4013_ (.Y(_1010_),
    .A(net948),
    .B(net376));
 sg13g2_and2_1 _4014_ (.A(net948),
    .B(net549),
    .X(_1011_));
 sg13g2_xor2_1 _4015_ (.B(net550),
    .A(net948),
    .X(_1012_));
 sg13g2_o21ai_1 _4016_ (.B1(_1007_),
    .Y(_1013_),
    .A1(_1005_),
    .A2(_1006_));
 sg13g2_xnor2_1 _4017_ (.Y(_1014_),
    .A(_1012_),
    .B(_1013_));
 sg13g2_o21ai_1 _4018_ (.B1(_1010_),
    .Y(_0060_),
    .A1(net372),
    .A2(_1014_));
 sg13g2_nand2_1 _4019_ (.Y(_1015_),
    .A(net961),
    .B(net377));
 sg13g2_a21oi_1 _4020_ (.A1(_1012_),
    .A2(_1013_),
    .Y(_1016_),
    .B1(_1011_));
 sg13g2_nor2_1 _4021_ (.A(net961),
    .B(net549),
    .Y(_1017_));
 sg13g2_nand2_1 _4022_ (.Y(_1018_),
    .A(net961),
    .B(net549));
 sg13g2_nand2b_1 _4023_ (.Y(_1019_),
    .B(_1018_),
    .A_N(_1017_));
 sg13g2_xnor2_1 _4024_ (.Y(_1020_),
    .A(_1016_),
    .B(_1019_));
 sg13g2_o21ai_1 _4025_ (.B1(_1015_),
    .Y(_0061_),
    .A1(net372),
    .A2(_1020_));
 sg13g2_nand2_1 _4026_ (.Y(_1021_),
    .A(net952),
    .B(net377));
 sg13g2_nor2b_1 _4027_ (.A(net549),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[6] ),
    .Y(_1022_));
 sg13g2_xnor2_1 _4028_ (.Y(_1023_),
    .A(net952),
    .B(net549));
 sg13g2_o21ai_1 _4029_ (.B1(_1018_),
    .Y(_1024_),
    .A1(_1016_),
    .A2(_1017_));
 sg13g2_xnor2_1 _4030_ (.Y(_1025_),
    .A(_1023_),
    .B(_1024_));
 sg13g2_o21ai_1 _4031_ (.B1(_1021_),
    .Y(_0062_),
    .A1(net373),
    .A2(_1025_));
 sg13g2_nand2_1 _4032_ (.Y(_1026_),
    .A(net885),
    .B(net376));
 sg13g2_a21oi_1 _4033_ (.A1(_1023_),
    .A2(_1024_),
    .Y(_1027_),
    .B1(_1022_));
 sg13g2_nand2b_1 _4034_ (.Y(_1028_),
    .B(net551),
    .A_N(net885));
 sg13g2_nand2_1 _4035_ (.Y(_1029_),
    .A(_0937_),
    .B(_1028_));
 sg13g2_xnor2_1 _4036_ (.Y(_1030_),
    .A(_1027_),
    .B(_1029_));
 sg13g2_o21ai_1 _4037_ (.B1(_1026_),
    .Y(_0063_),
    .A1(net373),
    .A2(_1030_));
 sg13g2_nand2_1 _4038_ (.Y(_1031_),
    .A(net918),
    .B(net376));
 sg13g2_nand2b_1 _4039_ (.Y(_1032_),
    .B(net548),
    .A_N(net918));
 sg13g2_nand2_1 _4040_ (.Y(_1033_),
    .A(_0937_),
    .B(_1027_));
 sg13g2_nand4_1 _4041_ (.B(_1028_),
    .C(_1032_),
    .A(_0939_),
    .Y(_1034_),
    .D(_1033_));
 sg13g2_a22oi_1 _4042_ (.Y(_1035_),
    .B1(_1033_),
    .B2(_1028_),
    .A2(_1032_),
    .A1(_0939_));
 sg13g2_nand2_1 _4043_ (.Y(_1036_),
    .A(_0992_),
    .B(_1034_));
 sg13g2_o21ai_1 _4044_ (.B1(_1031_),
    .Y(_0064_),
    .A1(_1035_),
    .A2(_1036_));
 sg13g2_nand2_1 _4045_ (.Y(_1037_),
    .A(_0939_),
    .B(_1034_));
 sg13g2_nand2b_1 _4046_ (.Y(_1038_),
    .B(net1012),
    .A_N(net548));
 sg13g2_nand2b_1 _4047_ (.Y(_1039_),
    .B(net548),
    .A_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[9] ));
 sg13g2_nand2_1 _4048_ (.Y(_1040_),
    .A(_1037_),
    .B(_1039_));
 sg13g2_nor2b_1 _4049_ (.A(_1040_),
    .B_N(_1038_),
    .Y(_1041_));
 sg13g2_a21oi_1 _4050_ (.A1(_1038_),
    .A2(_1039_),
    .Y(_1042_),
    .B1(_1037_));
 sg13g2_nor3_1 _4051_ (.A(net372),
    .B(_1041_),
    .C(_1042_),
    .Y(_1043_));
 sg13g2_a21o_1 _4052_ (.A2(net376),
    .A1(net1012),
    .B1(_1043_),
    .X(_0065_));
 sg13g2_nand2_1 _4053_ (.Y(_1044_),
    .A(net982),
    .B(net376));
 sg13g2_nand2_1 _4054_ (.Y(_1045_),
    .A(_1038_),
    .B(_1040_));
 sg13g2_or2_1 _4055_ (.X(_1046_),
    .B(net548),
    .A(net982));
 sg13g2_xnor2_1 _4056_ (.Y(_1047_),
    .A(net982),
    .B(net548));
 sg13g2_xnor2_1 _4057_ (.Y(_1048_),
    .A(_1045_),
    .B(_1047_));
 sg13g2_o21ai_1 _4058_ (.B1(_1044_),
    .Y(_0066_),
    .A1(net372),
    .A2(_1048_));
 sg13g2_nor2_1 _4059_ (.A(_0532_),
    .B(net423),
    .Y(_0082_));
 sg13g2_nand4_1 _4060_ (.B(net1012),
    .C(net548),
    .A(net982),
    .Y(_1049_),
    .D(_1037_));
 sg13g2_o21ai_1 _4061_ (.B1(_1049_),
    .Y(_1050_),
    .A1(_1045_),
    .A2(_1046_));
 sg13g2_a21oi_1 _4062_ (.A1(_0992_),
    .A2(_1050_),
    .Y(_1051_),
    .B1(_0082_));
 sg13g2_nand3_1 _4063_ (.B(_0987_),
    .C(_1050_),
    .A(net803),
    .Y(_1052_));
 sg13g2_nor2b_1 _4064_ (.A(_1051_),
    .B_N(_1052_),
    .Y(_0067_));
 sg13g2_and2_1 _4065_ (.A(net449),
    .B(net15),
    .X(_0068_));
 sg13g2_and2_1 _4066_ (.A(net449),
    .B(net16),
    .X(_0069_));
 sg13g2_nor2b_1 _4067_ (.A(net879),
    .B_N(_0987_),
    .Y(_1053_));
 sg13g2_mux2_1 _4068_ (.A0(_0992_),
    .A1(net378),
    .S(net879),
    .X(_0070_));
 sg13g2_nand2b_1 _4069_ (.Y(_1054_),
    .B(_1053_),
    .A_N(net840));
 sg13g2_xor2_1 _4070_ (.B(_1053_),
    .A(net840),
    .X(_1055_));
 sg13g2_and2_1 _4071_ (.A(net445),
    .B(_1055_),
    .X(_0071_));
 sg13g2_nand2_1 _4072_ (.Y(_1056_),
    .A(_0523_),
    .B(_1054_));
 sg13g2_or3_1 _4073_ (.A(net919),
    .B(net840),
    .C(net879),
    .X(_1057_));
 sg13g2_o21ai_1 _4074_ (.B1(_1056_),
    .Y(_0072_),
    .A1(net373),
    .A2(_1057_));
 sg13g2_nor2_1 _4075_ (.A(net919),
    .B(_1054_),
    .Y(_1058_));
 sg13g2_nor3_1 _4076_ (.A(net849),
    .B(net919),
    .C(_1054_),
    .Y(_1059_));
 sg13g2_xor2_1 _4077_ (.B(_1058_),
    .A(net849),
    .X(_1060_));
 sg13g2_and2_1 _4078_ (.A(net445),
    .B(_1060_),
    .X(_0073_));
 sg13g2_xor2_1 _4079_ (.B(_1059_),
    .A(net846),
    .X(_1061_));
 sg13g2_and2_1 _4080_ (.A(net445),
    .B(_1061_),
    .X(_0074_));
 sg13g2_or3_1 _4081_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[4] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[3] ),
    .C(_1057_),
    .X(_1062_));
 sg13g2_a21o_1 _4082_ (.A2(_1062_),
    .A1(_0987_),
    .B1(net824),
    .X(_1063_));
 sg13g2_nand3_1 _4083_ (.B(_0986_),
    .C(_1062_),
    .A(net824),
    .Y(_1064_));
 sg13g2_and3_1 _4084_ (.X(_0075_),
    .A(net445),
    .B(_1063_),
    .C(_1064_));
 sg13g2_and2_1 _4085_ (.A(_0531_),
    .B(_1064_),
    .X(_1065_));
 sg13g2_nor2_2 _4086_ (.A(_0531_),
    .B(_1064_),
    .Y(_1066_));
 sg13g2_nor3_1 _4087_ (.A(net420),
    .B(_1065_),
    .C(_1066_),
    .Y(_0076_));
 sg13g2_o21ai_1 _4088_ (.B1(net445),
    .Y(_1067_),
    .A1(net828),
    .A2(_1066_));
 sg13g2_a21oi_1 _4089_ (.A1(net828),
    .A2(_1066_),
    .Y(_0077_),
    .B1(_1067_));
 sg13g2_a21oi_1 _4090_ (.A1(net828),
    .A2(_1066_),
    .Y(_1068_),
    .B1(net821));
 sg13g2_and3_2 _4091_ (.X(_1069_),
    .A(net821),
    .B(net828),
    .C(_1066_));
 sg13g2_nor3_1 _4092_ (.A(net420),
    .B(_1068_),
    .C(_1069_),
    .Y(_0078_));
 sg13g2_xnor2_1 _4093_ (.Y(_1070_),
    .A(net865),
    .B(_1069_));
 sg13g2_nor2_1 _4094_ (.A(net419),
    .B(_1070_),
    .Y(_0079_));
 sg13g2_a21o_1 _4095_ (.A2(_1069_),
    .A1(net865),
    .B1(net859),
    .X(_1071_));
 sg13g2_nand3_1 _4096_ (.B(net865),
    .C(_1069_),
    .A(net859),
    .Y(_1072_));
 sg13g2_and3_1 _4097_ (.X(_0080_),
    .A(net441),
    .B(_1071_),
    .C(_1072_));
 sg13g2_xor2_1 _4098_ (.B(_1072_),
    .A(net878),
    .X(_1073_));
 sg13g2_nor2_1 _4099_ (.A(net419),
    .B(_1073_),
    .Y(_0081_));
 sg13g2_and2_1 _4100_ (.A(net498),
    .B(net798),
    .X(_0083_));
 sg13g2_nor2_1 _4101_ (.A(net799),
    .B(net435),
    .Y(_0084_));
 sg13g2_nor2b_1 _4102_ (.A(net532),
    .B_N(net834),
    .Y(_1074_));
 sg13g2_xnor2_1 _4103_ (.Y(_1075_),
    .A(net532),
    .B(net834));
 sg13g2_o21ai_1 _4104_ (.B1(net499),
    .Y(_1076_),
    .A1(net799),
    .A2(_1075_));
 sg13g2_a21oi_1 _4105_ (.A1(net799),
    .A2(_1075_),
    .Y(_0085_),
    .B1(_1076_));
 sg13g2_a21oi_1 _4106_ (.A1(net799),
    .A2(_1075_),
    .Y(_1077_),
    .B1(_1074_));
 sg13g2_nand2_1 _4107_ (.Y(_1078_),
    .A(net532),
    .B(net1057));
 sg13g2_xnor2_1 _4108_ (.Y(_1079_),
    .A(net532),
    .B(net1057));
 sg13g2_or2_1 _4109_ (.X(_1080_),
    .B(_1079_),
    .A(_1077_));
 sg13g2_nand2_1 _4110_ (.Y(_1081_),
    .A(net499),
    .B(_1080_));
 sg13g2_a21oi_1 _4111_ (.A1(_1077_),
    .A2(net1058),
    .Y(_0086_),
    .B1(_1081_));
 sg13g2_nand2_1 _4112_ (.Y(_1082_),
    .A(_0582_),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][4] ));
 sg13g2_xor2_1 _4113_ (.B(net1266),
    .A(net532),
    .X(_1083_));
 sg13g2_nand3_1 _4114_ (.B(_1080_),
    .C(_1083_),
    .A(_1078_),
    .Y(_1084_));
 sg13g2_a21o_1 _4115_ (.A2(_1080_),
    .A1(_1078_),
    .B1(_1083_),
    .X(_1085_));
 sg13g2_and3_1 _4116_ (.X(_0087_),
    .A(net499),
    .B(_1084_),
    .C(_1085_));
 sg13g2_and2_1 _4117_ (.A(_1082_),
    .B(_1085_),
    .X(_1086_));
 sg13g2_nand2_1 _4118_ (.Y(_1087_),
    .A(_0582_),
    .B(net1060));
 sg13g2_xor2_1 _4119_ (.B(net1060),
    .A(net533),
    .X(_1088_));
 sg13g2_or2_1 _4120_ (.X(_1089_),
    .B(_1088_),
    .A(_1086_));
 sg13g2_nand2_1 _4121_ (.Y(_1090_),
    .A(net501),
    .B(_1089_));
 sg13g2_a21oi_1 _4122_ (.A1(_1086_),
    .A2(_1088_),
    .Y(_0088_),
    .B1(_1090_));
 sg13g2_xor2_1 _4123_ (.B(net1222),
    .A(net533),
    .X(_1091_));
 sg13g2_a21oi_1 _4124_ (.A1(_1087_),
    .A2(_1089_),
    .Y(_1092_),
    .B1(_1091_));
 sg13g2_and3_1 _4125_ (.X(_1093_),
    .A(_1087_),
    .B(_1089_),
    .C(_1091_));
 sg13g2_nor3_1 _4126_ (.A(net436),
    .B(_1092_),
    .C(_1093_),
    .Y(_0089_));
 sg13g2_nor2_1 _4127_ (.A(_1089_),
    .B(_1091_),
    .Y(_1094_));
 sg13g2_o21ai_1 _4128_ (.B1(_1087_),
    .Y(_1095_),
    .A1(net533),
    .A2(_0589_));
 sg13g2_nor2_1 _4129_ (.A(_1094_),
    .B(_1095_),
    .Y(_1096_));
 sg13g2_nand2_1 _4130_ (.Y(_1097_),
    .A(_0582_),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][7] ));
 sg13g2_xor2_1 _4131_ (.B(net1175),
    .A(net533),
    .X(_1098_));
 sg13g2_or2_1 _4132_ (.X(_1099_),
    .B(_1098_),
    .A(_1096_));
 sg13g2_nand2_1 _4133_ (.Y(_1100_),
    .A(net501),
    .B(_1099_));
 sg13g2_a21oi_1 _4134_ (.A1(_1096_),
    .A2(_1098_),
    .Y(_0090_),
    .B1(_1100_));
 sg13g2_xor2_1 _4135_ (.B(net1149),
    .A(net534),
    .X(_1101_));
 sg13g2_and3_1 _4136_ (.X(_1102_),
    .A(_1097_),
    .B(_1099_),
    .C(_1101_));
 sg13g2_a21oi_1 _4137_ (.A1(_1097_),
    .A2(_1099_),
    .Y(_1103_),
    .B1(net1150));
 sg13g2_nor3_1 _4138_ (.A(net437),
    .B(_1102_),
    .C(net1151),
    .Y(_0091_));
 sg13g2_nor4_1 _4139_ (.A(_1089_),
    .B(_1091_),
    .C(_1098_),
    .D(_1101_),
    .Y(_1104_));
 sg13g2_o21ai_1 _4140_ (.B1(_1097_),
    .Y(_1105_),
    .A1(net533),
    .A2(_0590_));
 sg13g2_nor3_1 _4141_ (.A(_1095_),
    .B(_1104_),
    .C(_1105_),
    .Y(_1106_));
 sg13g2_xor2_1 _4142_ (.B(net1115),
    .A(net533),
    .X(_1107_));
 sg13g2_or2_1 _4143_ (.X(_1108_),
    .B(_1107_),
    .A(_1106_));
 sg13g2_nand2_1 _4144_ (.Y(_1109_),
    .A(net501),
    .B(_1108_));
 sg13g2_a21oi_1 _4145_ (.A1(_1106_),
    .A2(_1107_),
    .Y(_0092_),
    .B1(_1109_));
 sg13g2_o21ai_1 _4146_ (.B1(_1108_),
    .Y(_1110_),
    .A1(net533),
    .A2(_0591_));
 sg13g2_xnor2_1 _4147_ (.Y(_1111_),
    .A(net533),
    .B(net1036));
 sg13g2_o21ai_1 _4148_ (.B1(net501),
    .Y(_1112_),
    .A1(_1110_),
    .A2(_1111_));
 sg13g2_a21oi_1 _4149_ (.A1(_1110_),
    .A2(_1111_),
    .Y(_0093_),
    .B1(_1112_));
 sg13g2_nand2b_1 _4150_ (.Y(_1113_),
    .B(_1111_),
    .A_N(_1108_));
 sg13g2_o21ai_1 _4151_ (.B1(_0582_),
    .Y(_1114_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][9] ),
    .A2(net1036));
 sg13g2_and3_1 _4152_ (.X(_0094_),
    .A(net504),
    .B(_1113_),
    .C(net1037));
 sg13g2_nor2b_1 _4153_ (.A(net1103),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][6] ),
    .Y(_1115_));
 sg13g2_xnor2_1 _4154_ (.Y(_1116_),
    .A(net1103),
    .B(net1106));
 sg13g2_nor2_1 _4155_ (.A(net437),
    .B(_1116_),
    .Y(_0095_));
 sg13g2_nor2b_1 _4156_ (.A(net534),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][6] ),
    .Y(_1117_));
 sg13g2_xnor2_1 _4157_ (.Y(_1118_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][7] ),
    .B(_1117_));
 sg13g2_nand2_1 _4158_ (.Y(_1119_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][1] ),
    .B(_1118_));
 sg13g2_xnor2_1 _4159_ (.Y(_1120_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][1] ),
    .B(_1118_));
 sg13g2_o21ai_1 _4160_ (.B1(net495),
    .Y(_1121_),
    .A1(net1104),
    .A2(_1120_));
 sg13g2_a21oi_1 _4161_ (.A1(net1104),
    .A2(_1120_),
    .Y(_0096_),
    .B1(_1121_));
 sg13g2_o21ai_1 _4162_ (.B1(_1119_),
    .Y(_1122_),
    .A1(_1115_),
    .A2(_1120_));
 sg13g2_o21ai_1 _4163_ (.B1(_0582_),
    .Y(_1123_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][6] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][7] ));
 sg13g2_xnor2_1 _4164_ (.Y(_1124_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][8] ),
    .B(_1123_));
 sg13g2_nor2b_1 _4165_ (.A(_1124_),
    .B_N(net1355),
    .Y(_1125_));
 sg13g2_xnor2_1 _4166_ (.Y(_1126_),
    .A(net1355),
    .B(_1124_));
 sg13g2_nor2_1 _4167_ (.A(_1122_),
    .B(_1126_),
    .Y(_1127_));
 sg13g2_a21oi_1 _4168_ (.A1(_1122_),
    .A2(_1126_),
    .Y(_1128_),
    .B1(net439));
 sg13g2_nor2b_1 _4169_ (.A(net1356),
    .B_N(_1128_),
    .Y(_0097_));
 sg13g2_a21o_1 _4170_ (.A2(_1126_),
    .A1(_1122_),
    .B1(_1125_),
    .X(_1129_));
 sg13g2_o21ai_1 _4171_ (.B1(_1123_),
    .Y(_1130_),
    .A1(net534),
    .A2(_0586_));
 sg13g2_nor2b_1 _4172_ (.A(net534),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][9] ),
    .Y(_1131_));
 sg13g2_xnor2_1 _4173_ (.Y(_1132_),
    .A(net1574),
    .B(_1130_));
 sg13g2_and2_1 _4174_ (.A(net1363),
    .B(_1132_),
    .X(_1133_));
 sg13g2_xor2_1 _4175_ (.B(_1132_),
    .A(net1363),
    .X(_1134_));
 sg13g2_o21ai_1 _4176_ (.B1(net495),
    .Y(_1135_),
    .A1(_1129_),
    .A2(_1134_));
 sg13g2_a21oi_1 _4177_ (.A1(_1129_),
    .A2(net1364),
    .Y(_0098_),
    .B1(_1135_));
 sg13g2_a21o_1 _4178_ (.A2(_1134_),
    .A1(_1129_),
    .B1(_1133_),
    .X(_1136_));
 sg13g2_nor3_1 _4179_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][10] ),
    .B(_1130_),
    .C(_1131_),
    .Y(_1137_));
 sg13g2_o21ai_1 _4180_ (.B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][10] ),
    .Y(_1138_),
    .A1(_1130_),
    .A2(_1131_));
 sg13g2_nor2b_1 _4181_ (.A(_1137_),
    .B_N(_1138_),
    .Y(_1139_));
 sg13g2_nor2b_1 _4182_ (.A(_1139_),
    .B_N(net1499),
    .Y(_1140_));
 sg13g2_nand2b_1 _4183_ (.Y(_1141_),
    .B(_1139_),
    .A_N(net1499));
 sg13g2_nand2b_1 _4184_ (.Y(_1142_),
    .B(_1141_),
    .A_N(_1140_));
 sg13g2_nor2b_1 _4185_ (.A(_1136_),
    .B_N(_1142_),
    .Y(_1143_));
 sg13g2_nor2b_1 _4186_ (.A(_1142_),
    .B_N(_1136_),
    .Y(_1144_));
 sg13g2_nor3_1 _4187_ (.A(net437),
    .B(_1143_),
    .C(_1144_),
    .Y(_0099_));
 sg13g2_a21o_2 _4188_ (.A2(_1141_),
    .A1(_1136_),
    .B1(_1140_),
    .X(_1145_));
 sg13g2_nor2_1 _4189_ (.A(net534),
    .B(_1137_),
    .Y(_1146_));
 sg13g2_xnor2_1 _4190_ (.Y(_1147_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][11] ),
    .B(_1146_));
 sg13g2_and2_1 _4191_ (.A(net1398),
    .B(_1147_),
    .X(_1148_));
 sg13g2_xor2_1 _4192_ (.B(_1147_),
    .A(net1398),
    .X(_1149_));
 sg13g2_o21ai_1 _4193_ (.B1(net495),
    .Y(_1150_),
    .A1(_1145_),
    .A2(_1149_));
 sg13g2_a21oi_1 _4194_ (.A1(_1145_),
    .A2(_1149_),
    .Y(_0100_),
    .B1(_1150_));
 sg13g2_a21oi_2 _4195_ (.B1(_1148_),
    .Y(_1151_),
    .A2(_1149_),
    .A1(_1145_));
 sg13g2_a21oi_1 _4196_ (.A1(_0587_),
    .A2(_1137_),
    .Y(_1152_),
    .B1(net534));
 sg13g2_nor2b_1 _4197_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][12] ),
    .B_N(_1152_),
    .Y(_1153_));
 sg13g2_xnor2_1 _4198_ (.Y(_1154_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][12] ),
    .B(_1152_));
 sg13g2_nand2_1 _4199_ (.Y(_1155_),
    .A(net991),
    .B(_1154_));
 sg13g2_xnor2_1 _4200_ (.Y(_1156_),
    .A(net991),
    .B(_1154_));
 sg13g2_or2_1 _4201_ (.X(_1157_),
    .B(_1156_),
    .A(_1151_));
 sg13g2_nand2_1 _4202_ (.Y(_1158_),
    .A(net496),
    .B(_1157_));
 sg13g2_a21oi_1 _4203_ (.A1(_1151_),
    .A2(_1156_),
    .Y(_0101_),
    .B1(_1158_));
 sg13g2_a21oi_1 _4204_ (.A1(net531),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][12] ),
    .Y(_1159_),
    .B1(_1153_));
 sg13g2_nor2_1 _4205_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[1] ),
    .B(net382),
    .Y(_1160_));
 sg13g2_xnor2_1 _4206_ (.Y(_1161_),
    .A(net1208),
    .B(net382));
 sg13g2_and3_1 _4207_ (.X(_1162_),
    .A(_1155_),
    .B(_1157_),
    .C(_1161_));
 sg13g2_a21oi_1 _4208_ (.A1(_1155_),
    .A2(_1157_),
    .Y(_1163_),
    .B1(_1161_));
 sg13g2_nor3_1 _4209_ (.A(net433),
    .B(_1162_),
    .C(_1163_),
    .Y(_0102_));
 sg13g2_nor3_1 _4210_ (.A(_1151_),
    .B(_1156_),
    .C(_1160_),
    .Y(_1164_));
 sg13g2_a221oi_1 _4211_ (.B2(net1208),
    .C1(_1164_),
    .B1(net382),
    .A1(net991),
    .Y(_1165_),
    .A2(_1154_));
 sg13g2_xnor2_1 _4212_ (.Y(_1166_),
    .A(net1183),
    .B(net382));
 sg13g2_nor2_1 _4213_ (.A(_1165_),
    .B(_1166_),
    .Y(_1167_));
 sg13g2_a21oi_1 _4214_ (.A1(_1165_),
    .A2(_1166_),
    .Y(_1168_),
    .B1(net433));
 sg13g2_nor2b_1 _4215_ (.A(_1167_),
    .B_N(_1168_),
    .Y(_0103_));
 sg13g2_xnor2_1 _4216_ (.Y(_1169_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[3] ),
    .B(net382));
 sg13g2_a21oi_1 _4217_ (.A1(net1183),
    .A2(net382),
    .Y(_1170_),
    .B1(_1167_));
 sg13g2_o21ai_1 _4218_ (.B1(net486),
    .Y(_1171_),
    .A1(_1169_),
    .A2(_1170_));
 sg13g2_a21oi_1 _4219_ (.A1(_1169_),
    .A2(_1170_),
    .Y(_0104_),
    .B1(_1171_));
 sg13g2_xnor2_1 _4220_ (.Y(_1172_),
    .A(net1300),
    .B(net383));
 sg13g2_or3_1 _4221_ (.A(_1165_),
    .B(_1166_),
    .C(_1169_),
    .X(_1173_));
 sg13g2_o21ai_1 _4222_ (.B1(net383),
    .Y(_1174_),
    .A1(net1183),
    .A2(net1559));
 sg13g2_and2_1 _4223_ (.A(_1173_),
    .B(_1174_),
    .X(_1175_));
 sg13g2_and2_1 _4224_ (.A(_1172_),
    .B(_1175_),
    .X(_1176_));
 sg13g2_nor2_1 _4225_ (.A(_1172_),
    .B(_1175_),
    .Y(_1177_));
 sg13g2_nor3_1 _4226_ (.A(net433),
    .B(_1176_),
    .C(_1177_),
    .Y(_0105_));
 sg13g2_xnor2_1 _4227_ (.Y(_1178_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[5] ),
    .B(net383));
 sg13g2_a21oi_1 _4228_ (.A1(net1300),
    .A2(net382),
    .Y(_1179_),
    .B1(_1177_));
 sg13g2_o21ai_1 _4229_ (.B1(net496),
    .Y(_1180_),
    .A1(_1178_),
    .A2(_1179_));
 sg13g2_a21oi_1 _4230_ (.A1(_1178_),
    .A2(_1179_),
    .Y(_0106_),
    .B1(_1180_));
 sg13g2_nor3_1 _4231_ (.A(_1172_),
    .B(_1173_),
    .C(_1178_),
    .Y(_1181_));
 sg13g2_o21ai_1 _4232_ (.B1(net382),
    .Y(_1182_),
    .A1(net1300),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[5] ));
 sg13g2_nand2_1 _4233_ (.Y(_1183_),
    .A(_1174_),
    .B(_1182_));
 sg13g2_nor2_1 _4234_ (.A(_1181_),
    .B(_1183_),
    .Y(_1184_));
 sg13g2_xnor2_1 _4235_ (.Y(_1185_),
    .A(net1309),
    .B(net383));
 sg13g2_o21ai_1 _4236_ (.B1(net496),
    .Y(_1186_),
    .A1(_1184_),
    .A2(_1185_));
 sg13g2_a21oi_1 _4237_ (.A1(_1184_),
    .A2(_1185_),
    .Y(_0107_),
    .B1(_1186_));
 sg13g2_nand2_1 _4238_ (.Y(_1187_),
    .A(net962),
    .B(net991));
 sg13g2_o21ai_1 _4239_ (.B1(net479),
    .Y(_1188_),
    .A1(net962),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[0] ));
 sg13g2_nor2b_1 _4240_ (.A(net963),
    .B_N(_1187_),
    .Y(_0108_));
 sg13g2_nor2b_1 _4241_ (.A(net531),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[0] ),
    .Y(_1189_));
 sg13g2_xnor2_1 _4242_ (.Y(_1190_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[1] ),
    .B(_1189_));
 sg13g2_or2_1 _4243_ (.X(_1191_),
    .B(_1190_),
    .A(_0583_));
 sg13g2_xnor2_1 _4244_ (.Y(_1192_),
    .A(_0583_),
    .B(_1190_));
 sg13g2_o21ai_1 _4245_ (.B1(net479),
    .Y(_1193_),
    .A1(_1187_),
    .A2(_1192_));
 sg13g2_a21oi_1 _4246_ (.A1(_1187_),
    .A2(_1192_),
    .Y(_0109_),
    .B1(_1193_));
 sg13g2_o21ai_1 _4247_ (.B1(_1191_),
    .Y(_1194_),
    .A1(_1187_),
    .A2(_1192_));
 sg13g2_o21ai_1 _4248_ (.B1(_0582_),
    .Y(_1195_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[0] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[1] ));
 sg13g2_xnor2_1 _4249_ (.Y(_1196_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[2] ),
    .B(_1195_));
 sg13g2_and2_1 _4250_ (.A(net1277),
    .B(_1196_),
    .X(_1197_));
 sg13g2_xor2_1 _4251_ (.B(_1196_),
    .A(net1277),
    .X(_1198_));
 sg13g2_nor2_1 _4252_ (.A(_1194_),
    .B(net1278),
    .Y(_1199_));
 sg13g2_a21oi_1 _4253_ (.A1(_1194_),
    .A2(_1198_),
    .Y(_1200_),
    .B1(net429));
 sg13g2_nor2b_1 _4254_ (.A(net1279),
    .B_N(_1200_),
    .Y(_0110_));
 sg13g2_a21oi_1 _4255_ (.A1(_1194_),
    .A2(_1198_),
    .Y(_1201_),
    .B1(_1197_));
 sg13g2_o21ai_1 _4256_ (.B1(_1195_),
    .Y(_1202_),
    .A1(net531),
    .A2(_0584_));
 sg13g2_xor2_1 _4257_ (.B(_1202_),
    .A(net1576),
    .X(_1203_));
 sg13g2_nand2_1 _4258_ (.Y(_1204_),
    .A(net1322),
    .B(_1203_));
 sg13g2_xnor2_1 _4259_ (.Y(_1205_),
    .A(net1322),
    .B(_1203_));
 sg13g2_o21ai_1 _4260_ (.B1(net479),
    .Y(_1206_),
    .A1(_1201_),
    .A2(_1205_));
 sg13g2_a21oi_1 _4261_ (.A1(_1201_),
    .A2(_1205_),
    .Y(_0111_),
    .B1(_1206_));
 sg13g2_o21ai_1 _4262_ (.B1(_1204_),
    .Y(_1207_),
    .A1(_1201_),
    .A2(_1205_));
 sg13g2_nor2b_1 _4263_ (.A(net531),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[3] ),
    .Y(_1208_));
 sg13g2_nor2_1 _4264_ (.A(_1202_),
    .B(_1208_),
    .Y(_1209_));
 sg13g2_nor3_1 _4265_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[4] ),
    .B(_1202_),
    .C(_1208_),
    .Y(_1210_));
 sg13g2_xnor2_1 _4266_ (.Y(_1211_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[4] ),
    .B(_1209_));
 sg13g2_and2_1 _4267_ (.A(net1501),
    .B(_1211_),
    .X(_1212_));
 sg13g2_or2_1 _4268_ (.X(_1213_),
    .B(_1211_),
    .A(net1501));
 sg13g2_nor2b_1 _4269_ (.A(_1212_),
    .B_N(_1213_),
    .Y(_1214_));
 sg13g2_nor2_1 _4270_ (.A(_1207_),
    .B(_1214_),
    .Y(_1215_));
 sg13g2_a21oi_1 _4271_ (.A1(_1207_),
    .A2(_1214_),
    .Y(_1216_),
    .B1(net435));
 sg13g2_nor2b_1 _4272_ (.A(_1215_),
    .B_N(_1216_),
    .Y(_0112_));
 sg13g2_a21oi_1 _4273_ (.A1(_1207_),
    .A2(_1213_),
    .Y(_1217_),
    .B1(_1212_));
 sg13g2_nor2_1 _4274_ (.A(net531),
    .B(_1210_),
    .Y(_1218_));
 sg13g2_xnor2_1 _4275_ (.Y(_1219_),
    .A(_0585_),
    .B(_1218_));
 sg13g2_nand2_1 _4276_ (.Y(_1220_),
    .A(net1404),
    .B(_1219_));
 sg13g2_xnor2_1 _4277_ (.Y(_1221_),
    .A(net1404),
    .B(_1219_));
 sg13g2_o21ai_1 _4278_ (.B1(net497),
    .Y(_1222_),
    .A1(_1217_),
    .A2(_1221_));
 sg13g2_a21oi_1 _4279_ (.A1(_1217_),
    .A2(_1221_),
    .Y(_0113_),
    .B1(_1222_));
 sg13g2_o21ai_1 _4280_ (.B1(_1220_),
    .Y(_1223_),
    .A1(_1217_),
    .A2(_1221_));
 sg13g2_a21oi_1 _4281_ (.A1(_0585_),
    .A2(_1210_),
    .Y(_1224_),
    .B1(net531));
 sg13g2_nor2b_1 _4282_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[10] ),
    .B_N(_1224_),
    .Y(_1225_));
 sg13g2_xnor2_1 _4283_ (.Y(_1226_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[10] ),
    .B(_1224_));
 sg13g2_nor2b_1 _4284_ (.A(_1226_),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][6] ),
    .Y(_1227_));
 sg13g2_xor2_1 _4285_ (.B(_1226_),
    .A(net1106),
    .X(_1228_));
 sg13g2_inv_1 _4286_ (.Y(_1229_),
    .A(_1228_));
 sg13g2_nor2_1 _4287_ (.A(_1223_),
    .B(_1229_),
    .Y(_1230_));
 sg13g2_and2_1 _4288_ (.A(_1223_),
    .B(_1229_),
    .X(_1231_));
 sg13g2_nor3_1 _4289_ (.A(net435),
    .B(_1230_),
    .C(_1231_),
    .Y(_0114_));
 sg13g2_a21oi_1 _4290_ (.A1(_1223_),
    .A2(_1229_),
    .Y(_1232_),
    .B1(_1227_));
 sg13g2_a21oi_2 _4291_ (.B1(_1225_),
    .Y(_1233_),
    .A2(net1309),
    .A1(net531));
 sg13g2_inv_1 _4292_ (.Y(_1234_),
    .A(net381));
 sg13g2_nor2b_1 _4293_ (.A(net381),
    .B_N(net1567),
    .Y(_1235_));
 sg13g2_xnor2_1 _4294_ (.Y(_1236_),
    .A(net1462),
    .B(net381));
 sg13g2_nor2b_1 _4295_ (.A(_1236_),
    .B_N(_1232_),
    .Y(_1237_));
 sg13g2_nor2b_1 _4296_ (.A(_1232_),
    .B_N(_1236_),
    .Y(_1238_));
 sg13g2_nor3_1 _4297_ (.A(net437),
    .B(net1463),
    .C(_1238_),
    .Y(_0115_));
 sg13g2_xnor2_1 _4298_ (.Y(_1239_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][8] ),
    .B(net381));
 sg13g2_or3_1 _4299_ (.A(_1235_),
    .B(_1238_),
    .C(_1239_),
    .X(_1240_));
 sg13g2_o21ai_1 _4300_ (.B1(_1239_),
    .Y(_1241_),
    .A1(_1235_),
    .A2(_1238_));
 sg13g2_and3_1 _4301_ (.X(_0116_),
    .A(net501),
    .B(net1568),
    .C(_1241_));
 sg13g2_xor2_1 _4302_ (.B(net381),
    .A(net1512),
    .X(_1242_));
 sg13g2_inv_1 _4303_ (.Y(_1243_),
    .A(_1242_));
 sg13g2_o21ai_1 _4304_ (.B1(_1241_),
    .Y(_1244_),
    .A1(_0586_),
    .A2(net381));
 sg13g2_o21ai_1 _4305_ (.B1(net501),
    .Y(_1245_),
    .A1(_1243_),
    .A2(_1244_));
 sg13g2_a21oi_1 _4306_ (.A1(_1243_),
    .A2(_1244_),
    .Y(_0117_),
    .B1(_1245_));
 sg13g2_xnor2_1 _4307_ (.Y(_1246_),
    .A(net1527),
    .B(net381));
 sg13g2_nor2_1 _4308_ (.A(_1241_),
    .B(_1242_),
    .Y(_1247_));
 sg13g2_o21ai_1 _4309_ (.B1(_1234_),
    .Y(_1248_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][8] ),
    .A2(net1512));
 sg13g2_o21ai_1 _4310_ (.B1(_1248_),
    .Y(_1249_),
    .A1(_1241_),
    .A2(_1242_));
 sg13g2_nor2_1 _4311_ (.A(_1246_),
    .B(_1249_),
    .Y(_1250_));
 sg13g2_and2_1 _4312_ (.A(_1246_),
    .B(_1249_),
    .X(_1251_));
 sg13g2_nor3_1 _4313_ (.A(net437),
    .B(net1528),
    .C(_1251_),
    .Y(_0118_));
 sg13g2_xnor2_1 _4314_ (.Y(_1252_),
    .A(net1360),
    .B(_1233_));
 sg13g2_a21o_1 _4315_ (.A2(_1234_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][10] ),
    .B1(_1251_),
    .X(_1253_));
 sg13g2_o21ai_1 _4316_ (.B1(net501),
    .Y(_1254_),
    .A1(_1252_),
    .A2(_1253_));
 sg13g2_a21oi_1 _4317_ (.A1(net1361),
    .A2(_1253_),
    .Y(_0119_),
    .B1(_1254_));
 sg13g2_nand3_1 _4318_ (.B(_1247_),
    .C(_1252_),
    .A(_1246_),
    .Y(_1255_));
 sg13g2_o21ai_1 _4319_ (.B1(_1234_),
    .Y(_1256_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][10] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][11] ));
 sg13g2_nand3_1 _4320_ (.B(_1255_),
    .C(_1256_),
    .A(_1248_),
    .Y(_1257_));
 sg13g2_xnor2_1 _4321_ (.Y(_1258_),
    .A(net1199),
    .B(net381));
 sg13g2_o21ai_1 _4322_ (.B1(net497),
    .Y(_1259_),
    .A1(_1257_),
    .A2(_1258_));
 sg13g2_a21oi_1 _4323_ (.A1(_1257_),
    .A2(_1258_),
    .Y(_0120_),
    .B1(_1259_));
 sg13g2_nor2_1 _4324_ (.A(net770),
    .B(net436),
    .Y(_0121_));
 sg13g2_nor2b_1 _4325_ (.A(net542),
    .B_N(net817),
    .Y(_1260_));
 sg13g2_xnor2_1 _4326_ (.Y(_1261_),
    .A(net542),
    .B(net817));
 sg13g2_o21ai_1 _4327_ (.B1(net498),
    .Y(_1262_),
    .A1(net770),
    .A2(_1261_));
 sg13g2_a21oi_1 _4328_ (.A1(net770),
    .A2(_1261_),
    .Y(_0122_),
    .B1(_1262_));
 sg13g2_a21oi_1 _4329_ (.A1(net770),
    .A2(_1261_),
    .Y(_1263_),
    .B1(_1260_));
 sg13g2_nand2_1 _4330_ (.Y(_1264_),
    .A(net542),
    .B(net1026));
 sg13g2_xnor2_1 _4331_ (.Y(_1265_),
    .A(net542),
    .B(net1026));
 sg13g2_or2_1 _4332_ (.X(_1266_),
    .B(_1265_),
    .A(_1263_));
 sg13g2_nand2_1 _4333_ (.Y(_1267_),
    .A(net502),
    .B(_1266_));
 sg13g2_a21oi_1 _4334_ (.A1(_1263_),
    .A2(net1027),
    .Y(_0123_),
    .B1(_1267_));
 sg13g2_nand2_1 _4335_ (.Y(_1268_),
    .A(net410),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][3] ));
 sg13g2_xor2_1 _4336_ (.B(net1284),
    .A(net542),
    .X(_1269_));
 sg13g2_nand3_1 _4337_ (.B(_1266_),
    .C(_1269_),
    .A(_1264_),
    .Y(_1270_));
 sg13g2_a21o_1 _4338_ (.A2(_1266_),
    .A1(_1264_),
    .B1(_1269_),
    .X(_1271_));
 sg13g2_and3_1 _4339_ (.X(_0124_),
    .A(net502),
    .B(_1270_),
    .C(_1271_));
 sg13g2_and2_1 _4340_ (.A(_1268_),
    .B(_1271_),
    .X(_1272_));
 sg13g2_nand2_1 _4341_ (.Y(_1273_),
    .A(net410),
    .B(net1080));
 sg13g2_xor2_1 _4342_ (.B(net1080),
    .A(net541),
    .X(_1274_));
 sg13g2_or2_1 _4343_ (.X(_1275_),
    .B(_1274_),
    .A(_1272_));
 sg13g2_nand2_1 _4344_ (.Y(_1276_),
    .A(net502),
    .B(_1275_));
 sg13g2_a21oi_1 _4345_ (.A1(_1272_),
    .A2(_1274_),
    .Y(_0125_),
    .B1(_1276_));
 sg13g2_xor2_1 _4346_ (.B(net1120),
    .A(net541),
    .X(_1277_));
 sg13g2_a21oi_1 _4347_ (.A1(_1273_),
    .A2(_1275_),
    .Y(_1278_),
    .B1(_1277_));
 sg13g2_and3_1 _4348_ (.X(_1279_),
    .A(_1273_),
    .B(_1275_),
    .C(_1277_));
 sg13g2_nor3_1 _4349_ (.A(net436),
    .B(_1278_),
    .C(_1279_),
    .Y(_0126_));
 sg13g2_nor2_1 _4350_ (.A(_1275_),
    .B(_1277_),
    .Y(_1280_));
 sg13g2_o21ai_1 _4351_ (.B1(_1273_),
    .Y(_1281_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].z_sign ),
    .A2(_0606_));
 sg13g2_nor2_1 _4352_ (.A(_1280_),
    .B(_1281_),
    .Y(_1282_));
 sg13g2_nand2_1 _4353_ (.Y(_1283_),
    .A(net410),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][6] ));
 sg13g2_xor2_1 _4354_ (.B(net1192),
    .A(net541),
    .X(_1284_));
 sg13g2_or2_1 _4355_ (.X(_1285_),
    .B(_1284_),
    .A(_1282_));
 sg13g2_nand2_1 _4356_ (.Y(_1286_),
    .A(net503),
    .B(_1285_));
 sg13g2_a21oi_1 _4357_ (.A1(_1282_),
    .A2(_1284_),
    .Y(_0127_),
    .B1(_1286_));
 sg13g2_xor2_1 _4358_ (.B(net1138),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].z_sign ),
    .X(_1287_));
 sg13g2_and3_1 _4359_ (.X(_1288_),
    .A(_1283_),
    .B(_1285_),
    .C(_1287_));
 sg13g2_a21oi_1 _4360_ (.A1(_1283_),
    .A2(_1285_),
    .Y(_1289_),
    .B1(net1139));
 sg13g2_nor3_1 _4361_ (.A(net436),
    .B(_1288_),
    .C(net1140),
    .Y(_0128_));
 sg13g2_nor2_1 _4362_ (.A(_1284_),
    .B(_1287_),
    .Y(_1290_));
 sg13g2_nand2b_1 _4363_ (.Y(_1291_),
    .B(_1283_),
    .A_N(_1281_));
 sg13g2_a221oi_1 _4364_ (.B2(_1290_),
    .C1(_1291_),
    .B1(_1280_),
    .A1(net411),
    .Y(_1292_),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][7] ));
 sg13g2_xor2_1 _4365_ (.B(net1110),
    .A(net541),
    .X(_1293_));
 sg13g2_or2_1 _4366_ (.X(_1294_),
    .B(_1293_),
    .A(_1292_));
 sg13g2_nand2_1 _4367_ (.Y(_1295_),
    .A(net503),
    .B(_1294_));
 sg13g2_a21oi_1 _4368_ (.A1(_1292_),
    .A2(_1293_),
    .Y(_0129_),
    .B1(_1295_));
 sg13g2_o21ai_1 _4369_ (.B1(_1294_),
    .Y(_1296_),
    .A1(net541),
    .A2(_0607_));
 sg13g2_xnor2_1 _4370_ (.Y(_1297_),
    .A(net541),
    .B(net1121));
 sg13g2_o21ai_1 _4371_ (.B1(net503),
    .Y(_1298_),
    .A1(_1296_),
    .A2(_1297_));
 sg13g2_a21oi_1 _4372_ (.A1(_1296_),
    .A2(_1297_),
    .Y(_0130_),
    .B1(_1298_));
 sg13g2_nand2b_1 _4373_ (.Y(_1299_),
    .B(_1297_),
    .A_N(_1294_));
 sg13g2_o21ai_1 _4374_ (.B1(net410),
    .Y(_1300_),
    .A1(net1110),
    .A2(net1121));
 sg13g2_and2_1 _4375_ (.A(_1299_),
    .B(_1300_),
    .X(_1301_));
 sg13g2_xor2_1 _4376_ (.B(net818),
    .A(net541),
    .X(_1302_));
 sg13g2_o21ai_1 _4377_ (.B1(net501),
    .Y(_1303_),
    .A1(_1301_),
    .A2(_1302_));
 sg13g2_a21oi_1 _4378_ (.A1(_1301_),
    .A2(_1302_),
    .Y(_0131_),
    .B1(_1303_));
 sg13g2_a21oi_1 _4379_ (.A1(net410),
    .A2(net818),
    .Y(_0132_),
    .B1(_1303_));
 sg13g2_nor2b_1 _4380_ (.A(net922),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][7] ),
    .Y(_1304_));
 sg13g2_xnor2_1 _4381_ (.Y(_1305_),
    .A(net922),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][7] ));
 sg13g2_nor2_1 _4382_ (.A(net435),
    .B(net923),
    .Y(_0133_));
 sg13g2_nor2b_1 _4383_ (.A(net542),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][7] ),
    .Y(_1306_));
 sg13g2_xnor2_1 _4384_ (.Y(_1307_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][8] ),
    .B(_1306_));
 sg13g2_nand2_1 _4385_ (.Y(_1308_),
    .A(net1097),
    .B(_1307_));
 sg13g2_xnor2_1 _4386_ (.Y(_1309_),
    .A(net1097),
    .B(_1307_));
 sg13g2_o21ai_1 _4387_ (.B1(net502),
    .Y(_1310_),
    .A1(_1304_),
    .A2(_1309_));
 sg13g2_a21oi_1 _4388_ (.A1(_1304_),
    .A2(_1309_),
    .Y(_0134_),
    .B1(_1310_));
 sg13g2_o21ai_1 _4389_ (.B1(_1308_),
    .Y(_1311_),
    .A1(_1304_),
    .A2(_1309_));
 sg13g2_or2_1 _4390_ (.X(_1312_),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][8] ),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][7] ));
 sg13g2_a21o_1 _4391_ (.A2(_1312_),
    .A1(net410),
    .B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][9] ),
    .X(_1313_));
 sg13g2_nand3_1 _4392_ (.B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][9] ),
    .C(_1312_),
    .A(net410),
    .Y(_1314_));
 sg13g2_a21oi_1 _4393_ (.A1(_1313_),
    .A2(_1314_),
    .Y(_1315_),
    .B1(_0604_));
 sg13g2_nand3_1 _4394_ (.B(_1313_),
    .C(_1314_),
    .A(_0604_),
    .Y(_1316_));
 sg13g2_nor2b_1 _4395_ (.A(_1315_),
    .B_N(_1316_),
    .Y(_1317_));
 sg13g2_nor2_1 _4396_ (.A(_1311_),
    .B(_1317_),
    .Y(_1318_));
 sg13g2_a21oi_1 _4397_ (.A1(_1311_),
    .A2(_1317_),
    .Y(_1319_),
    .B1(net436));
 sg13g2_nor2b_1 _4398_ (.A(_1318_),
    .B_N(_1319_),
    .Y(_0135_));
 sg13g2_a21o_1 _4399_ (.A2(_1317_),
    .A1(_1311_),
    .B1(_1315_),
    .X(_1320_));
 sg13g2_o21ai_1 _4400_ (.B1(net410),
    .Y(_1321_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][9] ),
    .A2(_1312_));
 sg13g2_xnor2_1 _4401_ (.Y(_1322_),
    .A(_0603_),
    .B(_1321_));
 sg13g2_and2_1 _4402_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][3] ),
    .B(_1322_),
    .X(_1323_));
 sg13g2_xor2_1 _4403_ (.B(_1322_),
    .A(net1452),
    .X(_1324_));
 sg13g2_o21ai_1 _4404_ (.B1(net497),
    .Y(_1325_),
    .A1(_1320_),
    .A2(_1324_));
 sg13g2_a21oi_1 _4405_ (.A1(_1320_),
    .A2(_1324_),
    .Y(_0136_),
    .B1(_1325_));
 sg13g2_a21o_1 _4406_ (.A2(_1324_),
    .A1(_1320_),
    .B1(_1323_),
    .X(_1326_));
 sg13g2_o21ai_1 _4407_ (.B1(_1321_),
    .Y(_1327_),
    .A1(net542),
    .A2(_0603_));
 sg13g2_nor2_1 _4408_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][11] ),
    .B(_1327_),
    .Y(_1328_));
 sg13g2_xnor2_1 _4409_ (.Y(_1329_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][11] ),
    .B(_1327_));
 sg13g2_and2_1 _4410_ (.A(net1374),
    .B(_1329_),
    .X(_1330_));
 sg13g2_xor2_1 _4411_ (.B(_1329_),
    .A(net1374),
    .X(_1331_));
 sg13g2_nor2_1 _4412_ (.A(_1326_),
    .B(_1331_),
    .Y(_1332_));
 sg13g2_a21oi_1 _4413_ (.A1(_1326_),
    .A2(_1331_),
    .Y(_1333_),
    .B1(net435));
 sg13g2_nor2b_1 _4414_ (.A(net1375),
    .B_N(_1333_),
    .Y(_0137_));
 sg13g2_a21oi_1 _4415_ (.A1(_1326_),
    .A2(_1331_),
    .Y(_1334_),
    .B1(_1330_));
 sg13g2_nor3_1 _4416_ (.A(net543),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][12] ),
    .C(_1328_),
    .Y(_1335_));
 sg13g2_o21ai_1 _4417_ (.B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][12] ),
    .Y(_1336_),
    .A1(net543),
    .A2(_1328_));
 sg13g2_nor2b_1 _4418_ (.A(_1335_),
    .B_N(_1336_),
    .Y(_1337_));
 sg13g2_nand2_1 _4419_ (.Y(_1338_),
    .A(net1411),
    .B(_1337_));
 sg13g2_xnor2_1 _4420_ (.Y(_1339_),
    .A(net1411),
    .B(_1337_));
 sg13g2_or2_1 _4421_ (.X(_1340_),
    .B(_1339_),
    .A(_1334_));
 sg13g2_nand2_1 _4422_ (.Y(_1341_),
    .A(net496),
    .B(_1340_));
 sg13g2_a21oi_1 _4423_ (.A1(_1334_),
    .A2(_1339_),
    .Y(_0138_),
    .B1(_1341_));
 sg13g2_a21oi_1 _4424_ (.A1(net543),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][12] ),
    .Y(_1342_),
    .B1(_1335_));
 sg13g2_and2_1 _4425_ (.A(net1471),
    .B(net387),
    .X(_1343_));
 sg13g2_xnor2_1 _4426_ (.Y(_1344_),
    .A(net1471),
    .B(net387));
 sg13g2_and3_1 _4427_ (.X(_1345_),
    .A(_1338_),
    .B(_1340_),
    .C(_1344_));
 sg13g2_a21oi_1 _4428_ (.A1(_1338_),
    .A2(_1340_),
    .Y(_1346_),
    .B1(_1344_));
 sg13g2_a21o_1 _4429_ (.A2(_1340_),
    .A1(_1338_),
    .B1(_1344_),
    .X(_1347_));
 sg13g2_nor3_1 _4430_ (.A(net433),
    .B(_1345_),
    .C(_1346_),
    .Y(_0139_));
 sg13g2_nand2b_1 _4431_ (.Y(_1348_),
    .B(_1347_),
    .A_N(_1343_));
 sg13g2_nand2_1 _4432_ (.Y(_1349_),
    .A(net996),
    .B(net386));
 sg13g2_or2_1 _4433_ (.X(_1350_),
    .B(net387),
    .A(net996));
 sg13g2_and2_1 _4434_ (.A(_1349_),
    .B(_1350_),
    .X(_1351_));
 sg13g2_o21ai_1 _4435_ (.B1(net487),
    .Y(_1352_),
    .A1(_1348_),
    .A2(_1351_));
 sg13g2_a21oi_1 _4436_ (.A1(_1348_),
    .A2(_1351_),
    .Y(_0140_),
    .B1(_1352_));
 sg13g2_nand2_1 _4437_ (.Y(_1353_),
    .A(net1472),
    .B(net386));
 sg13g2_xnor2_1 _4438_ (.Y(_1354_),
    .A(net1472),
    .B(net386));
 sg13g2_o21ai_1 _4439_ (.B1(_1350_),
    .Y(_1355_),
    .A1(_1343_),
    .A2(_1346_));
 sg13g2_nand3_1 _4440_ (.B(_1354_),
    .C(_1355_),
    .A(_1349_),
    .Y(_1356_));
 sg13g2_a21o_1 _4441_ (.A2(_1355_),
    .A1(_1349_),
    .B1(_1354_),
    .X(_1357_));
 sg13g2_and3_1 _4442_ (.X(_0141_),
    .A(net486),
    .B(_1356_),
    .C(_1357_));
 sg13g2_xnor2_1 _4443_ (.Y(_1358_),
    .A(net1369),
    .B(net386));
 sg13g2_and2_1 _4444_ (.A(_1353_),
    .B(_1357_),
    .X(_1359_));
 sg13g2_o21ai_1 _4445_ (.B1(net486),
    .Y(_1360_),
    .A1(_1358_),
    .A2(_1359_));
 sg13g2_a21oi_1 _4446_ (.A1(_1358_),
    .A2(_1359_),
    .Y(_0142_),
    .B1(_1360_));
 sg13g2_nor2_1 _4447_ (.A(_1357_),
    .B(_1358_),
    .Y(_1361_));
 sg13g2_o21ai_1 _4448_ (.B1(net386),
    .Y(_1362_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[1] ),
    .A2(net1369));
 sg13g2_nor2b_1 _4449_ (.A(_1361_),
    .B_N(net1370),
    .Y(_1363_));
 sg13g2_o21ai_1 _4450_ (.B1(_1362_),
    .Y(_1364_),
    .A1(_1357_),
    .A2(_1358_));
 sg13g2_xnor2_1 _4451_ (.Y(_1365_),
    .A(net1158),
    .B(net386));
 sg13g2_nor2b_1 _4452_ (.A(_1365_),
    .B_N(_1364_),
    .Y(_1366_));
 sg13g2_nand2b_1 _4453_ (.Y(_1367_),
    .B(net486),
    .A_N(_1366_));
 sg13g2_a21oi_1 _4454_ (.A1(_1363_),
    .A2(_1365_),
    .Y(_0143_),
    .B1(_1367_));
 sg13g2_xnor2_1 _4455_ (.Y(_1368_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[4] ),
    .B(net386));
 sg13g2_a21oi_1 _4456_ (.A1(net1158),
    .A2(net386),
    .Y(_1369_),
    .B1(_1366_));
 sg13g2_o21ai_1 _4457_ (.B1(net486),
    .Y(_1370_),
    .A1(_1368_),
    .A2(_1369_));
 sg13g2_a21oi_1 _4458_ (.A1(_1368_),
    .A2(_1369_),
    .Y(_0144_),
    .B1(_1370_));
 sg13g2_nor2_1 _4459_ (.A(_1365_),
    .B(_1368_),
    .Y(_1371_));
 sg13g2_o21ai_1 _4460_ (.B1(net387),
    .Y(_1372_),
    .A1(net1158),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[4] ));
 sg13g2_nand2_1 _4461_ (.Y(_1373_),
    .A(_1362_),
    .B(_1372_));
 sg13g2_a21oi_1 _4462_ (.A1(_1361_),
    .A2(_1371_),
    .Y(_1374_),
    .B1(_1373_));
 sg13g2_xnor2_1 _4463_ (.Y(_1375_),
    .A(net1287),
    .B(net387));
 sg13g2_o21ai_1 _4464_ (.B1(net486),
    .Y(_1376_),
    .A1(_1374_),
    .A2(_1375_));
 sg13g2_a21oi_1 _4465_ (.A1(_1374_),
    .A2(_1375_),
    .Y(_0145_),
    .B1(_1376_));
 sg13g2_nand2_1 _4466_ (.Y(_1377_),
    .A(net985),
    .B(net996));
 sg13g2_o21ai_1 _4467_ (.B1(net486),
    .Y(_1378_),
    .A1(net985),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[0] ));
 sg13g2_nor2b_1 _4468_ (.A(net986),
    .B_N(_1377_),
    .Y(_0146_));
 sg13g2_nand2b_1 _4469_ (.Y(_1379_),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[0] ),
    .A_N(net543));
 sg13g2_xnor2_1 _4470_ (.Y(_1380_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[1] ),
    .B(_1379_));
 sg13g2_nand2_1 _4471_ (.Y(_1381_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][1] ),
    .B(_1380_));
 sg13g2_xnor2_1 _4472_ (.Y(_1382_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][1] ),
    .B(_1380_));
 sg13g2_o21ai_1 _4473_ (.B1(net487),
    .Y(_1383_),
    .A1(_1377_),
    .A2(_1382_));
 sg13g2_a21oi_1 _4474_ (.A1(_1377_),
    .A2(_1382_),
    .Y(_0147_),
    .B1(_1383_));
 sg13g2_o21ai_1 _4475_ (.B1(_1381_),
    .Y(_1384_),
    .A1(_1377_),
    .A2(_1382_));
 sg13g2_or2_1 _4476_ (.X(_1385_),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[1] ),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[0] ));
 sg13g2_nand2_1 _4477_ (.Y(_1386_),
    .A(net411),
    .B(_1385_));
 sg13g2_a21oi_1 _4478_ (.A1(net411),
    .A2(_1385_),
    .Y(_1387_),
    .B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[2] ));
 sg13g2_xnor2_1 _4479_ (.Y(_1388_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[2] ),
    .B(_1386_));
 sg13g2_and2_1 _4480_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][2] ),
    .B(_1388_),
    .X(_1389_));
 sg13g2_xor2_1 _4481_ (.B(_1388_),
    .A(net1223),
    .X(_1390_));
 sg13g2_nor2_1 _4482_ (.A(_1384_),
    .B(net1224),
    .Y(_1391_));
 sg13g2_a21oi_1 _4483_ (.A1(_1384_),
    .A2(_1390_),
    .Y(_1392_),
    .B1(net433));
 sg13g2_nor2b_1 _4484_ (.A(net1225),
    .B_N(_1392_),
    .Y(_0148_));
 sg13g2_a21oi_1 _4485_ (.A1(_1384_),
    .A2(_1390_),
    .Y(_1393_),
    .B1(_1389_));
 sg13g2_nor2_1 _4486_ (.A(net543),
    .B(_1387_),
    .Y(_1394_));
 sg13g2_xnor2_1 _4487_ (.Y(_1395_),
    .A(_0601_),
    .B(_1394_));
 sg13g2_nand2_1 _4488_ (.Y(_1396_),
    .A(net1206),
    .B(_1395_));
 sg13g2_xnor2_1 _4489_ (.Y(_1397_),
    .A(net1206),
    .B(_1395_));
 sg13g2_or2_1 _4490_ (.X(_1398_),
    .B(_1397_),
    .A(_1393_));
 sg13g2_nand2_1 _4491_ (.Y(_1399_),
    .A(net486),
    .B(_1398_));
 sg13g2_a21oi_1 _4492_ (.A1(_1393_),
    .A2(_1397_),
    .Y(_0149_),
    .B1(_1399_));
 sg13g2_and2_1 _4493_ (.A(_1396_),
    .B(_1398_),
    .X(_1400_));
 sg13g2_o21ai_1 _4494_ (.B1(_1396_),
    .Y(_1401_),
    .A1(_1393_),
    .A2(_1397_));
 sg13g2_a21oi_1 _4495_ (.A1(_0601_),
    .A2(_1387_),
    .Y(_1402_),
    .B1(net543));
 sg13g2_nor2_1 _4496_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[4] ),
    .B(_1402_),
    .Y(_1403_));
 sg13g2_xnor2_1 _4497_ (.Y(_1404_),
    .A(net1480),
    .B(_1402_));
 sg13g2_nor2_1 _4498_ (.A(_0602_),
    .B(_1404_),
    .Y(_1405_));
 sg13g2_nand2_1 _4499_ (.Y(_1406_),
    .A(_0602_),
    .B(_1404_));
 sg13g2_nand2b_1 _4500_ (.Y(_1407_),
    .B(net1442),
    .A_N(_1405_));
 sg13g2_o21ai_1 _4501_ (.B1(net489),
    .Y(_1408_),
    .A1(_1400_),
    .A2(_1407_));
 sg13g2_a21oi_1 _4502_ (.A1(_1400_),
    .A2(_1407_),
    .Y(_0150_),
    .B1(_1408_));
 sg13g2_a21oi_1 _4503_ (.A1(_1401_),
    .A2(_1406_),
    .Y(_1409_),
    .B1(_1405_));
 sg13g2_nor2_1 _4504_ (.A(net543),
    .B(_1403_),
    .Y(_1410_));
 sg13g2_xnor2_1 _4505_ (.Y(_1411_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[10] ),
    .B(_1410_));
 sg13g2_nand2b_1 _4506_ (.Y(_1412_),
    .B(net1461),
    .A_N(_1411_));
 sg13g2_xor2_1 _4507_ (.B(_1411_),
    .A(net1461),
    .X(_1413_));
 sg13g2_o21ai_1 _4508_ (.B1(net498),
    .Y(_1414_),
    .A1(_1409_),
    .A2(_1413_));
 sg13g2_a21oi_1 _4509_ (.A1(_1409_),
    .A2(_1413_),
    .Y(_0151_),
    .B1(_1414_));
 sg13g2_o21ai_1 _4510_ (.B1(_1412_),
    .Y(_1415_),
    .A1(_1409_),
    .A2(_1413_));
 sg13g2_mux2_1 _4511_ (.A0(_1410_),
    .A1(net543),
    .S(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[10] ),
    .X(_1416_));
 sg13g2_and2_1 _4512_ (.A(net1332),
    .B(net384),
    .X(_1417_));
 sg13g2_xor2_1 _4513_ (.B(net384),
    .A(net1332),
    .X(_1418_));
 sg13g2_nor2_1 _4514_ (.A(_1415_),
    .B(_1418_),
    .Y(_1419_));
 sg13g2_a21oi_1 _4515_ (.A1(_1415_),
    .A2(_1418_),
    .Y(_1420_),
    .B1(net438));
 sg13g2_nor2b_1 _4516_ (.A(_1419_),
    .B_N(_1420_),
    .Y(_0152_));
 sg13g2_a21oi_1 _4517_ (.A1(_1415_),
    .A2(_1418_),
    .Y(_1421_),
    .B1(_1417_));
 sg13g2_nor2_1 _4518_ (.A(net1537),
    .B(net384),
    .Y(_1422_));
 sg13g2_xnor2_1 _4519_ (.Y(_1423_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][7] ),
    .B(net384));
 sg13g2_o21ai_1 _4520_ (.B1(net498),
    .Y(_1424_),
    .A1(_1421_),
    .A2(_1423_));
 sg13g2_a21oi_1 _4521_ (.A1(_1421_),
    .A2(_1423_),
    .Y(_0153_),
    .B1(_1424_));
 sg13g2_xor2_1 _4522_ (.B(net384),
    .A(net1477),
    .X(_1425_));
 sg13g2_a221oi_1 _4523_ (.B2(_1415_),
    .C1(_1417_),
    .B1(_1418_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][7] ),
    .Y(_1426_),
    .A2(net384));
 sg13g2_nor2_1 _4524_ (.A(_1422_),
    .B(_1426_),
    .Y(_1427_));
 sg13g2_and2_1 _4525_ (.A(_1425_),
    .B(_1427_),
    .X(_1428_));
 sg13g2_o21ai_1 _4526_ (.B1(net498),
    .Y(_1429_),
    .A1(_1425_),
    .A2(_1427_));
 sg13g2_nor2_1 _4527_ (.A(_1428_),
    .B(_1429_),
    .Y(_0154_));
 sg13g2_xor2_1 _4528_ (.B(net385),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][9] ),
    .X(_1430_));
 sg13g2_a21o_1 _4529_ (.A2(net384),
    .A1(net1477),
    .B1(_1428_),
    .X(_1431_));
 sg13g2_o21ai_1 _4530_ (.B1(net499),
    .Y(_1432_),
    .A1(_1430_),
    .A2(_1431_));
 sg13g2_a21oi_1 _4531_ (.A1(_1430_),
    .A2(_1431_),
    .Y(_0155_),
    .B1(_1432_));
 sg13g2_nand2_1 _4532_ (.Y(_1433_),
    .A(_1428_),
    .B(_1430_));
 sg13g2_o21ai_1 _4533_ (.B1(net385),
    .Y(_1434_),
    .A1(net1477),
    .A2(net1532));
 sg13g2_xnor2_1 _4534_ (.Y(_1435_),
    .A(net1169),
    .B(net385));
 sg13g2_and3_1 _4535_ (.X(_1436_),
    .A(_1433_),
    .B(_1434_),
    .C(_1435_));
 sg13g2_a21oi_1 _4536_ (.A1(_1433_),
    .A2(_1434_),
    .Y(_1437_),
    .B1(_1435_));
 sg13g2_nor3_1 _4537_ (.A(net438),
    .B(_1436_),
    .C(_1437_),
    .Y(_0156_));
 sg13g2_xor2_1 _4538_ (.B(net385),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][11] ),
    .X(_1438_));
 sg13g2_inv_1 _4539_ (.Y(_1439_),
    .A(_1438_));
 sg13g2_a21oi_1 _4540_ (.A1(net1169),
    .A2(net384),
    .Y(_1440_),
    .B1(_1437_));
 sg13g2_o21ai_1 _4541_ (.B1(net498),
    .Y(_1441_),
    .A1(_1439_),
    .A2(_1440_));
 sg13g2_a21oi_1 _4542_ (.A1(_1439_),
    .A2(_1440_),
    .Y(_0157_),
    .B1(_1441_));
 sg13g2_or3_1 _4543_ (.A(_1433_),
    .B(_1435_),
    .C(_1439_),
    .X(_1442_));
 sg13g2_o21ai_1 _4544_ (.B1(net385),
    .Y(_1443_),
    .A1(net1169),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][11] ));
 sg13g2_and3_1 _4545_ (.X(_1444_),
    .A(_1434_),
    .B(_1442_),
    .C(_1443_));
 sg13g2_xnor2_1 _4546_ (.Y(_1445_),
    .A(net1262),
    .B(net385));
 sg13g2_o21ai_1 _4547_ (.B1(net498),
    .Y(_1446_),
    .A1(_1444_),
    .A2(_1445_));
 sg13g2_a21oi_1 _4548_ (.A1(_1444_),
    .A2(_1445_),
    .Y(_0158_),
    .B1(_1446_));
 sg13g2_nor2_1 _4549_ (.A(net760),
    .B(net436),
    .Y(_0159_));
 sg13g2_nand2_1 _4550_ (.Y(_1447_),
    .A(net539),
    .B(net1006));
 sg13g2_xor2_1 _4551_ (.B(net1006),
    .A(net539),
    .X(_1448_));
 sg13g2_nand2_1 _4552_ (.Y(_1449_),
    .A(net760),
    .B(_1448_));
 sg13g2_o21ai_1 _4553_ (.B1(net502),
    .Y(_1450_),
    .A1(net760),
    .A2(_1448_));
 sg13g2_nor2b_1 _4554_ (.A(_1450_),
    .B_N(_1449_),
    .Y(_0160_));
 sg13g2_xor2_1 _4555_ (.B(net1272),
    .A(net539),
    .X(_1451_));
 sg13g2_nand3_1 _4556_ (.B(_1449_),
    .C(_1451_),
    .A(_1447_),
    .Y(_1452_));
 sg13g2_a21o_1 _4557_ (.A2(_1449_),
    .A1(_1447_),
    .B1(_1451_),
    .X(_1453_));
 sg13g2_and3_1 _4558_ (.X(_0161_),
    .A(net502),
    .B(_1452_),
    .C(_1453_));
 sg13g2_o21ai_1 _4559_ (.B1(_1453_),
    .Y(_1454_),
    .A1(net539),
    .A2(_0611_));
 sg13g2_nor2b_1 _4560_ (.A(net539),
    .B_N(net1419),
    .Y(_1455_));
 sg13g2_nand2b_1 _4561_ (.Y(_1456_),
    .B(net539),
    .A_N(net1419));
 sg13g2_nor2b_1 _4562_ (.A(_1455_),
    .B_N(_1456_),
    .Y(_1457_));
 sg13g2_o21ai_1 _4563_ (.B1(net502),
    .Y(_1458_),
    .A1(_1454_),
    .A2(_1457_));
 sg13g2_a21oi_1 _4564_ (.A1(_1454_),
    .A2(_1457_),
    .Y(_0162_),
    .B1(_1458_));
 sg13g2_nand2_1 _4565_ (.Y(_1459_),
    .A(_0608_),
    .B(net1038));
 sg13g2_xor2_1 _4566_ (.B(net1038),
    .A(net539),
    .X(_1460_));
 sg13g2_o21ai_1 _4567_ (.B1(_1456_),
    .Y(_1461_),
    .A1(_1454_),
    .A2(_1455_));
 sg13g2_or2_1 _4568_ (.X(_1462_),
    .B(_1461_),
    .A(_1460_));
 sg13g2_nand2_1 _4569_ (.Y(_1463_),
    .A(net503),
    .B(_1462_));
 sg13g2_a21oi_1 _4570_ (.A1(_1460_),
    .A2(_1461_),
    .Y(_0163_),
    .B1(_1463_));
 sg13g2_xor2_1 _4571_ (.B(net1153),
    .A(net539),
    .X(_1464_));
 sg13g2_a21oi_1 _4572_ (.A1(_1459_),
    .A2(_1462_),
    .Y(_1465_),
    .B1(_1464_));
 sg13g2_and3_1 _4573_ (.X(_1466_),
    .A(_1459_),
    .B(_1462_),
    .C(_1464_));
 sg13g2_nor3_1 _4574_ (.A(net436),
    .B(_1465_),
    .C(_1466_),
    .Y(_0164_));
 sg13g2_nor2_1 _4575_ (.A(_1462_),
    .B(_1464_),
    .Y(_1467_));
 sg13g2_o21ai_1 _4576_ (.B1(_1459_),
    .Y(_1468_),
    .A1(net540),
    .A2(_0612_));
 sg13g2_nor2_1 _4577_ (.A(_1467_),
    .B(_1468_),
    .Y(_1469_));
 sg13g2_nand2_1 _4578_ (.Y(_1470_),
    .A(_0608_),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][6] ));
 sg13g2_xor2_1 _4579_ (.B(net1214),
    .A(net540),
    .X(_1471_));
 sg13g2_or2_1 _4580_ (.X(_1472_),
    .B(_1471_),
    .A(_1469_));
 sg13g2_nand2_1 _4581_ (.Y(_1473_),
    .A(net503),
    .B(_1472_));
 sg13g2_a21oi_1 _4582_ (.A1(_1469_),
    .A2(_1471_),
    .Y(_0165_),
    .B1(_1473_));
 sg13g2_xor2_1 _4583_ (.B(net1133),
    .A(net540),
    .X(_1474_));
 sg13g2_and3_1 _4584_ (.X(_1475_),
    .A(_1470_),
    .B(_1472_),
    .C(_1474_));
 sg13g2_a21oi_1 _4585_ (.A1(_1470_),
    .A2(_1472_),
    .Y(_1476_),
    .B1(net1134));
 sg13g2_nor3_1 _4586_ (.A(net437),
    .B(_1475_),
    .C(net1135),
    .Y(_0166_));
 sg13g2_nor2_1 _4587_ (.A(_1471_),
    .B(_1474_),
    .Y(_1477_));
 sg13g2_nand2b_1 _4588_ (.Y(_1478_),
    .B(_1470_),
    .A_N(_1468_));
 sg13g2_a221oi_1 _4589_ (.B2(_1477_),
    .C1(_1478_),
    .B1(_1467_),
    .A1(_0608_),
    .Y(_1479_),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][7] ));
 sg13g2_nand2_1 _4590_ (.Y(_1480_),
    .A(_0608_),
    .B(net1086));
 sg13g2_xor2_1 _4591_ (.B(net1086),
    .A(net540),
    .X(_1481_));
 sg13g2_or2_1 _4592_ (.X(_1482_),
    .B(_1481_),
    .A(_1479_));
 sg13g2_nand2_1 _4593_ (.Y(_1483_),
    .A(net503),
    .B(_1482_));
 sg13g2_a21oi_1 _4594_ (.A1(_1479_),
    .A2(net1087),
    .Y(_0167_),
    .B1(_1483_));
 sg13g2_xor2_1 _4595_ (.B(net1185),
    .A(net540),
    .X(_1484_));
 sg13g2_a21oi_1 _4596_ (.A1(_1480_),
    .A2(_1482_),
    .Y(_1485_),
    .B1(_1484_));
 sg13g2_and3_1 _4597_ (.X(_1486_),
    .A(_1480_),
    .B(_1482_),
    .C(_1484_));
 sg13g2_nor3_1 _4598_ (.A(net437),
    .B(_1485_),
    .C(_1486_),
    .Y(_0168_));
 sg13g2_o21ai_1 _4599_ (.B1(_1480_),
    .Y(_1487_),
    .A1(_1482_),
    .A2(_1484_));
 sg13g2_a21oi_1 _4600_ (.A1(_0608_),
    .A2(net1185),
    .Y(_1488_),
    .B1(_1487_));
 sg13g2_xor2_1 _4601_ (.B(net832),
    .A(net540),
    .X(_1489_));
 sg13g2_o21ai_1 _4602_ (.B1(net502),
    .Y(_1490_),
    .A1(_1488_),
    .A2(_1489_));
 sg13g2_a21oi_1 _4603_ (.A1(_1488_),
    .A2(_1489_),
    .Y(_0169_),
    .B1(_1490_));
 sg13g2_a21oi_1 _4604_ (.A1(_0608_),
    .A2(net832),
    .Y(_0170_),
    .B1(_1490_));
 sg13g2_nor2b_1 _4605_ (.A(net976),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][8] ),
    .Y(_1491_));
 sg13g2_xnor2_1 _4606_ (.Y(_1492_),
    .A(net976),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][8] ));
 sg13g2_nor2_1 _4607_ (.A(net438),
    .B(net977),
    .Y(_0171_));
 sg13g2_nor2b_1 _4608_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].z_sign ),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][8] ),
    .Y(_1493_));
 sg13g2_xnor2_1 _4609_ (.Y(_1494_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][9] ),
    .B(_1493_));
 sg13g2_nand2_1 _4610_ (.Y(_1495_),
    .A(net1165),
    .B(_1494_));
 sg13g2_xnor2_1 _4611_ (.Y(_1496_),
    .A(net1165),
    .B(_1494_));
 sg13g2_o21ai_1 _4612_ (.B1(net498),
    .Y(_1497_),
    .A1(_1491_),
    .A2(_1496_));
 sg13g2_a21oi_1 _4613_ (.A1(_1491_),
    .A2(_1496_),
    .Y(_0172_),
    .B1(_1497_));
 sg13g2_o21ai_1 _4614_ (.B1(_1495_),
    .Y(_1498_),
    .A1(_1491_),
    .A2(_1496_));
 sg13g2_nor2_1 _4615_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][8] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][9] ),
    .Y(_1499_));
 sg13g2_nor2_1 _4616_ (.A(net538),
    .B(_1499_),
    .Y(_1500_));
 sg13g2_xnor2_1 _4617_ (.Y(_1501_),
    .A(net1273),
    .B(_1500_));
 sg13g2_and2_1 _4618_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][2] ),
    .B(_1501_),
    .X(_1502_));
 sg13g2_xor2_1 _4619_ (.B(_1501_),
    .A(net1382),
    .X(_1503_));
 sg13g2_nor2_1 _4620_ (.A(_1498_),
    .B(_1503_),
    .Y(_1504_));
 sg13g2_a21oi_1 _4621_ (.A1(_1498_),
    .A2(_1503_),
    .Y(_1505_),
    .B1(net433));
 sg13g2_nor2b_1 _4622_ (.A(_1504_),
    .B_N(_1505_),
    .Y(_0173_));
 sg13g2_a21oi_1 _4623_ (.A1(_1498_),
    .A2(_1503_),
    .Y(_1506_),
    .B1(_1502_));
 sg13g2_nor3_1 _4624_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][8] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][9] ),
    .C(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][10] ),
    .Y(_1507_));
 sg13g2_nor2_1 _4625_ (.A(net538),
    .B(_1507_),
    .Y(_1508_));
 sg13g2_xnor2_1 _4626_ (.Y(_1509_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][11] ),
    .B(_1508_));
 sg13g2_xor2_1 _4627_ (.B(_1509_),
    .A(net1350),
    .X(_1510_));
 sg13g2_nor2b_1 _4628_ (.A(net1351),
    .B_N(_1506_),
    .Y(_1511_));
 sg13g2_nor2b_1 _4629_ (.A(_1506_),
    .B_N(_1510_),
    .Y(_1512_));
 sg13g2_nor3_1 _4630_ (.A(net433),
    .B(net1352),
    .C(_1512_),
    .Y(_0174_));
 sg13g2_a21oi_1 _4631_ (.A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][3] ),
    .A2(_1509_),
    .Y(_1513_),
    .B1(_1512_));
 sg13g2_nor2b_1 _4632_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][11] ),
    .B_N(_1507_),
    .Y(_1514_));
 sg13g2_nor3_1 _4633_ (.A(net537),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][12] ),
    .C(_1514_),
    .Y(_1515_));
 sg13g2_o21ai_1 _4634_ (.B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][12] ),
    .Y(_1516_),
    .A1(net537),
    .A2(_1514_));
 sg13g2_nor2b_2 _4635_ (.A(_1515_),
    .B_N(_1516_),
    .Y(_1517_));
 sg13g2_nand2_2 _4636_ (.Y(_1518_),
    .A(net1212),
    .B(_1517_));
 sg13g2_xnor2_1 _4637_ (.Y(_1519_),
    .A(net1212),
    .B(_1517_));
 sg13g2_or2_1 _4638_ (.X(_1520_),
    .B(_1519_),
    .A(_1513_));
 sg13g2_nand2_1 _4639_ (.Y(_1521_),
    .A(net481),
    .B(_1520_));
 sg13g2_a21oi_1 _4640_ (.A1(_1513_),
    .A2(_1519_),
    .Y(_0175_),
    .B1(_1521_));
 sg13g2_a21oi_1 _4641_ (.A1(net537),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][12] ),
    .Y(_1522_),
    .B1(_1515_));
 sg13g2_a21o_1 _4642_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][12] ),
    .A1(net537),
    .B1(_1515_),
    .X(_1523_));
 sg13g2_nand2_1 _4643_ (.Y(_1524_),
    .A(net1550),
    .B(net393));
 sg13g2_xnor2_1 _4644_ (.Y(_1525_),
    .A(net1271),
    .B(net393));
 sg13g2_a21oi_1 _4645_ (.A1(_1518_),
    .A2(_1520_),
    .Y(_1526_),
    .B1(_1525_));
 sg13g2_and3_1 _4646_ (.X(_1527_),
    .A(_1518_),
    .B(_1520_),
    .C(_1525_));
 sg13g2_nor3_1 _4647_ (.A(net432),
    .B(_1526_),
    .C(_1527_),
    .Y(_0176_));
 sg13g2_nand2_1 _4648_ (.Y(_1528_),
    .A(_1518_),
    .B(_1524_));
 sg13g2_nor2_1 _4649_ (.A(_1520_),
    .B(_1525_),
    .Y(_1529_));
 sg13g2_nor2_1 _4650_ (.A(_1528_),
    .B(_1529_),
    .Y(_1530_));
 sg13g2_nand2_1 _4651_ (.Y(_1531_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][6] ),
    .B(net393));
 sg13g2_xnor2_1 _4652_ (.Y(_1532_),
    .A(net1253),
    .B(net394));
 sg13g2_or2_1 _4653_ (.X(_1533_),
    .B(_1532_),
    .A(_1530_));
 sg13g2_nand2_1 _4654_ (.Y(_1534_),
    .A(net481),
    .B(_1533_));
 sg13g2_a21oi_1 _4655_ (.A1(_1530_),
    .A2(_1532_),
    .Y(_0177_),
    .B1(_1534_));
 sg13g2_xnor2_1 _4656_ (.Y(_1535_),
    .A(net1189),
    .B(net393));
 sg13g2_and3_1 _4657_ (.X(_1536_),
    .A(_1531_),
    .B(_1533_),
    .C(_1535_));
 sg13g2_a21oi_1 _4658_ (.A1(_1531_),
    .A2(_1533_),
    .Y(_1537_),
    .B1(_1535_));
 sg13g2_nor3_1 _4659_ (.A(net432),
    .B(_1536_),
    .C(net1190),
    .Y(_0178_));
 sg13g2_a21oi_1 _4660_ (.A1(_0610_),
    .A2(_1523_),
    .Y(_1538_),
    .B1(_1532_));
 sg13g2_nand3_1 _4661_ (.B(_1524_),
    .C(_1531_),
    .A(_1518_),
    .Y(_1539_));
 sg13g2_a221oi_1 _4662_ (.B2(_1538_),
    .C1(_1539_),
    .B1(_1529_),
    .A1(net1189),
    .Y(_1540_),
    .A2(net393));
 sg13g2_xnor2_1 _4663_ (.Y(_1541_),
    .A(net1017),
    .B(net393));
 sg13g2_and2_1 _4664_ (.A(_1540_),
    .B(_1541_),
    .X(_1542_));
 sg13g2_nor2_1 _4665_ (.A(_1540_),
    .B(_1541_),
    .Y(_1543_));
 sg13g2_nor3_1 _4666_ (.A(net432),
    .B(_1542_),
    .C(_1543_),
    .Y(_0179_));
 sg13g2_a21oi_1 _4667_ (.A1(net1017),
    .A2(net393),
    .Y(_1544_),
    .B1(_1543_));
 sg13g2_xnor2_1 _4668_ (.Y(_1545_),
    .A(net1188),
    .B(net394));
 sg13g2_o21ai_1 _4669_ (.B1(net485),
    .Y(_1546_),
    .A1(_1544_),
    .A2(_1545_));
 sg13g2_a21oi_1 _4670_ (.A1(_1544_),
    .A2(_1545_),
    .Y(_0180_),
    .B1(_1546_));
 sg13g2_xnor2_1 _4671_ (.Y(_1547_),
    .A(net1534),
    .B(net393));
 sg13g2_nand2b_1 _4672_ (.Y(_1548_),
    .B(_1543_),
    .A_N(_1545_));
 sg13g2_nor2_1 _4673_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[0] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[1] ),
    .Y(_1549_));
 sg13g2_nand2b_1 _4674_ (.Y(_1550_),
    .B(net394),
    .A_N(_1549_));
 sg13g2_and3_1 _4675_ (.X(_1551_),
    .A(_1547_),
    .B(_1548_),
    .C(_1550_));
 sg13g2_a21oi_1 _4676_ (.A1(_1548_),
    .A2(_1550_),
    .Y(_1552_),
    .B1(_1547_));
 sg13g2_nor3_1 _4677_ (.A(net432),
    .B(_1551_),
    .C(net1535),
    .Y(_0181_));
 sg13g2_a21oi_1 _4678_ (.A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[2] ),
    .A2(net394),
    .Y(_1553_),
    .B1(_1552_));
 sg13g2_and2_1 _4679_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[3] ),
    .B(_1523_),
    .X(_1554_));
 sg13g2_xnor2_1 _4680_ (.Y(_1555_),
    .A(net1177),
    .B(net394));
 sg13g2_o21ai_1 _4681_ (.B1(net485),
    .Y(_1556_),
    .A1(_1553_),
    .A2(_1555_));
 sg13g2_a21oi_1 _4682_ (.A1(_1553_),
    .A2(_1555_),
    .Y(_0182_),
    .B1(_1556_));
 sg13g2_nor2_1 _4683_ (.A(_1547_),
    .B(_1548_),
    .Y(_1557_));
 sg13g2_nor4_1 _4684_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[0] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[1] ),
    .C(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[2] ),
    .D(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[3] ),
    .Y(_1558_));
 sg13g2_and2_1 _4685_ (.A(net394),
    .B(_1558_),
    .X(_1559_));
 sg13g2_mux2_1 _4686_ (.A0(_1559_),
    .A1(_1554_),
    .S(_1557_),
    .X(_1560_));
 sg13g2_o21ai_1 _4687_ (.B1(net488),
    .Y(_1561_),
    .A1(net872),
    .A2(_1560_));
 sg13g2_a21oi_1 _4688_ (.A1(net872),
    .A2(_1560_),
    .Y(_0183_),
    .B1(_1561_));
 sg13g2_nand2_1 _4689_ (.Y(_1562_),
    .A(net993),
    .B(net1017));
 sg13g2_o21ai_1 _4690_ (.B1(net482),
    .Y(_1563_),
    .A1(net993),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[0] ));
 sg13g2_nor2b_1 _4691_ (.A(net994),
    .B_N(_1562_),
    .Y(_0184_));
 sg13g2_nand2b_1 _4692_ (.Y(_1564_),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[0] ),
    .A_N(net537));
 sg13g2_xnor2_1 _4693_ (.Y(_1565_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[1] ),
    .B(_1564_));
 sg13g2_nand2_1 _4694_ (.Y(_1566_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][1] ),
    .B(_1565_));
 sg13g2_xnor2_1 _4695_ (.Y(_1567_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][1] ),
    .B(_1565_));
 sg13g2_o21ai_1 _4696_ (.B1(net482),
    .Y(_1568_),
    .A1(_1562_),
    .A2(_1567_));
 sg13g2_a21oi_1 _4697_ (.A1(_1562_),
    .A2(_1567_),
    .Y(_0185_),
    .B1(_1568_));
 sg13g2_o21ai_1 _4698_ (.B1(_1566_),
    .Y(_1569_),
    .A1(_1562_),
    .A2(_1567_));
 sg13g2_nor2_1 _4699_ (.A(net537),
    .B(_1549_),
    .Y(_1570_));
 sg13g2_xnor2_1 _4700_ (.Y(_1571_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[2] ),
    .B(_1570_));
 sg13g2_nor2b_1 _4701_ (.A(_1571_),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][2] ),
    .Y(_1572_));
 sg13g2_xnor2_1 _4702_ (.Y(_1573_),
    .A(net1438),
    .B(_1571_));
 sg13g2_nor2_1 _4703_ (.A(_1569_),
    .B(_1573_),
    .Y(_1574_));
 sg13g2_a21oi_1 _4704_ (.A1(_1569_),
    .A2(_1573_),
    .Y(_1575_),
    .B1(net432));
 sg13g2_nor2b_1 _4705_ (.A(net1439),
    .B_N(_1575_),
    .Y(_0186_));
 sg13g2_a21oi_1 _4706_ (.A1(_1569_),
    .A2(_1573_),
    .Y(_1576_),
    .B1(_1572_));
 sg13g2_a21oi_1 _4707_ (.A1(_0609_),
    .A2(_1549_),
    .Y(_1577_),
    .B1(net537));
 sg13g2_xnor2_1 _4708_ (.Y(_1578_),
    .A(net1177),
    .B(_1577_));
 sg13g2_nand2b_1 _4709_ (.Y(_1579_),
    .B(net1311),
    .A_N(_1578_));
 sg13g2_xnor2_1 _4710_ (.Y(_1580_),
    .A(net1311),
    .B(_1578_));
 sg13g2_inv_1 _4711_ (.Y(_1581_),
    .A(_1580_));
 sg13g2_o21ai_1 _4712_ (.B1(net488),
    .Y(_1582_),
    .A1(_1576_),
    .A2(_1581_));
 sg13g2_a21oi_1 _4713_ (.A1(_1576_),
    .A2(_1581_),
    .Y(_0187_),
    .B1(_1582_));
 sg13g2_o21ai_1 _4714_ (.B1(_1579_),
    .Y(_1583_),
    .A1(_1576_),
    .A2(_1581_));
 sg13g2_nor2_1 _4715_ (.A(net537),
    .B(_1558_),
    .Y(_1584_));
 sg13g2_xnor2_1 _4716_ (.Y(_1585_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[10] ),
    .B(_1584_));
 sg13g2_nand2b_1 _4717_ (.Y(_1586_),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][4] ),
    .A_N(_1585_));
 sg13g2_inv_1 _4718_ (.Y(_1587_),
    .A(_1586_));
 sg13g2_xnor2_1 _4719_ (.Y(_1588_),
    .A(net1524),
    .B(_1585_));
 sg13g2_or2_1 _4720_ (.X(_1589_),
    .B(_1588_),
    .A(_1583_));
 sg13g2_nand2_1 _4721_ (.Y(_1590_),
    .A(_1583_),
    .B(_1588_));
 sg13g2_and3_1 _4722_ (.X(_0188_),
    .A(net488),
    .B(_1589_),
    .C(_1590_));
 sg13g2_nand2_1 _4723_ (.Y(_1591_),
    .A(_1586_),
    .B(_1590_));
 sg13g2_mux2_1 _4724_ (.A0(_1584_),
    .A1(net538),
    .S(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[10] ),
    .X(_1592_));
 sg13g2_nor2_1 _4725_ (.A(net1293),
    .B(net401),
    .Y(_1593_));
 sg13g2_xor2_1 _4726_ (.B(net401),
    .A(net1293),
    .X(_1594_));
 sg13g2_o21ai_1 _4727_ (.B1(net488),
    .Y(_1595_),
    .A1(_1591_),
    .A2(_1594_));
 sg13g2_a21oi_1 _4728_ (.A1(_1591_),
    .A2(_1594_),
    .Y(_0189_),
    .B1(_1595_));
 sg13g2_and2_1 _4729_ (.A(net1495),
    .B(net400),
    .X(_1596_));
 sg13g2_xnor2_1 _4730_ (.Y(_1597_),
    .A(net1495),
    .B(net400));
 sg13g2_a221oi_1 _4731_ (.B2(net1293),
    .C1(_1587_),
    .B1(net401),
    .A1(_1583_),
    .Y(_1598_),
    .A2(_1588_));
 sg13g2_o21ai_1 _4732_ (.B1(_1597_),
    .Y(_1599_),
    .A1(_1593_),
    .A2(_1598_));
 sg13g2_nor3_1 _4733_ (.A(_1593_),
    .B(_1597_),
    .C(_1598_),
    .Y(_1600_));
 sg13g2_nand2_1 _4734_ (.Y(_1601_),
    .A(net488),
    .B(net1496));
 sg13g2_nor2_1 _4735_ (.A(_1600_),
    .B(_1601_),
    .Y(_0190_));
 sg13g2_nor2_1 _4736_ (.A(_1596_),
    .B(_1600_),
    .Y(_1602_));
 sg13g2_nand2_1 _4737_ (.Y(_1603_),
    .A(net1458),
    .B(net400));
 sg13g2_or2_1 _4738_ (.X(_1604_),
    .B(net400),
    .A(net1458));
 sg13g2_nand2_1 _4739_ (.Y(_1605_),
    .A(_1603_),
    .B(_1604_));
 sg13g2_o21ai_1 _4740_ (.B1(net488),
    .Y(_1606_),
    .A1(_1602_),
    .A2(_1605_));
 sg13g2_a21oi_1 _4741_ (.A1(_1602_),
    .A2(_1605_),
    .Y(_0191_),
    .B1(_1606_));
 sg13g2_xnor2_1 _4742_ (.Y(_1607_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][8] ),
    .B(_1592_));
 sg13g2_o21ai_1 _4743_ (.B1(_1604_),
    .Y(_1608_),
    .A1(_1596_),
    .A2(_1600_));
 sg13g2_nand3_1 _4744_ (.B(_1607_),
    .C(_1608_),
    .A(_1603_),
    .Y(_1609_));
 sg13g2_a21oi_1 _4745_ (.A1(_1603_),
    .A2(_1608_),
    .Y(_1610_),
    .B1(_1607_));
 sg13g2_nand2_1 _4746_ (.Y(_1611_),
    .A(net489),
    .B(net1459));
 sg13g2_nor2_1 _4747_ (.A(_1610_),
    .B(_1611_),
    .Y(_0192_));
 sg13g2_a21o_1 _4748_ (.A2(net400),
    .A1(net1526),
    .B1(_1610_),
    .X(_1612_));
 sg13g2_xor2_1 _4749_ (.B(net401),
    .A(net1504),
    .X(_1613_));
 sg13g2_o21ai_1 _4750_ (.B1(net489),
    .Y(_1614_),
    .A1(_1612_),
    .A2(_1613_));
 sg13g2_a21oi_1 _4751_ (.A1(_1612_),
    .A2(_1613_),
    .Y(_0193_),
    .B1(_1614_));
 sg13g2_xor2_1 _4752_ (.B(net400),
    .A(net1273),
    .X(_1615_));
 sg13g2_nand2_1 _4753_ (.Y(_1616_),
    .A(_1610_),
    .B(_1613_));
 sg13g2_nand2b_1 _4754_ (.Y(_1617_),
    .B(net401),
    .A_N(_1499_));
 sg13g2_nand2_1 _4755_ (.Y(_1618_),
    .A(_1616_),
    .B(_1617_));
 sg13g2_nor2_1 _4756_ (.A(_1615_),
    .B(_1618_),
    .Y(_1619_));
 sg13g2_and2_1 _4757_ (.A(_1615_),
    .B(_1618_),
    .X(_1620_));
 sg13g2_nor3_1 _4758_ (.A(net433),
    .B(_1619_),
    .C(_1620_),
    .Y(_0194_));
 sg13g2_a21o_1 _4759_ (.A2(net400),
    .A1(net1273),
    .B1(_1620_),
    .X(_1621_));
 sg13g2_xor2_1 _4760_ (.B(net400),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][11] ),
    .X(_1622_));
 sg13g2_o21ai_1 _4761_ (.B1(net488),
    .Y(_1623_),
    .A1(_1621_),
    .A2(_1622_));
 sg13g2_a21oi_1 _4762_ (.A1(_1621_),
    .A2(_1622_),
    .Y(_0195_),
    .B1(_1623_));
 sg13g2_nand2_1 _4763_ (.Y(_1624_),
    .A(_1615_),
    .B(_1622_));
 sg13g2_nand2b_1 _4764_ (.Y(_1625_),
    .B(net401),
    .A_N(_1514_));
 sg13g2_o21ai_1 _4765_ (.B1(_1625_),
    .Y(_1626_),
    .A1(_1616_),
    .A2(_1624_));
 sg13g2_xor2_1 _4766_ (.B(net401),
    .A(net1399),
    .X(_1627_));
 sg13g2_o21ai_1 _4767_ (.B1(net488),
    .Y(_1628_),
    .A1(_1626_),
    .A2(_1627_));
 sg13g2_a21oi_1 _4768_ (.A1(_1626_),
    .A2(_1627_),
    .Y(_0196_),
    .B1(_1628_));
 sg13g2_nand4_1 _4769_ (.B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][2] ),
    .C(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][1] ),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][3] ),
    .Y(_1629_),
    .D(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][0] ));
 sg13g2_and4_1 _4770_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][7] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][6] ),
    .C(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][5] ),
    .D(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][4] ),
    .X(_1630_));
 sg13g2_nand3_1 _4771_ (.B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][8] ),
    .C(_1630_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][9] ),
    .Y(_1631_));
 sg13g2_o21ai_1 _4772_ (.B1(net536),
    .Y(_1632_),
    .A1(_1629_),
    .A2(_1631_));
 sg13g2_nor4_1 _4773_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][3] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][2] ),
    .C(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][1] ),
    .D(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][0] ),
    .Y(_1633_));
 sg13g2_nor2_1 _4774_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][9] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][8] ),
    .Y(_1634_));
 sg13g2_nor4_1 _4775_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][7] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][6] ),
    .C(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][5] ),
    .D(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][4] ),
    .Y(_1635_));
 sg13g2_nand3_1 _4776_ (.B(_1634_),
    .C(_1635_),
    .A(_1633_),
    .Y(_1636_));
 sg13g2_a221oi_1 _4777_ (.B2(_0613_),
    .C1(net436),
    .B1(_1636_),
    .A1(net1142),
    .Y(_0197_),
    .A2(_1632_));
 sg13g2_nor2b_1 _4778_ (.A(net1082),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][9] ),
    .Y(_1637_));
 sg13g2_xnor2_1 _4779_ (.Y(_1638_),
    .A(net1082),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][9] ));
 sg13g2_nor2_2 _4780_ (.A(net432),
    .B(net1083),
    .Y(_0198_));
 sg13g2_nor2b_1 _4781_ (.A(net536),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][9] ),
    .Y(_1639_));
 sg13g2_xnor2_1 _4782_ (.Y(_1640_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][10] ),
    .B(_1639_));
 sg13g2_nand2_1 _4783_ (.Y(_1641_),
    .A(net1365),
    .B(_1640_));
 sg13g2_xnor2_1 _4784_ (.Y(_1642_),
    .A(net1365),
    .B(_1640_));
 sg13g2_o21ai_1 _4785_ (.B1(net485),
    .Y(_1643_),
    .A1(_1637_),
    .A2(_1642_));
 sg13g2_a21oi_1 _4786_ (.A1(_1637_),
    .A2(_1642_),
    .Y(_0199_),
    .B1(_1643_));
 sg13g2_o21ai_1 _4787_ (.B1(_1641_),
    .Y(_1644_),
    .A1(_1637_),
    .A2(_1642_));
 sg13g2_or2_1 _4788_ (.X(_1645_),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][10] ),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][9] ));
 sg13g2_a21oi_1 _4789_ (.A1(_0613_),
    .A2(_1645_),
    .Y(_1646_),
    .B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][11] ));
 sg13g2_nand3_1 _4790_ (.B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][11] ),
    .C(_1645_),
    .A(_0613_),
    .Y(_1647_));
 sg13g2_nor2b_1 _4791_ (.A(_1646_),
    .B_N(_1647_),
    .Y(_1648_));
 sg13g2_nand2b_1 _4792_ (.Y(_1649_),
    .B(net1470),
    .A_N(_1648_));
 sg13g2_xnor2_1 _4793_ (.Y(_1650_),
    .A(net1470),
    .B(_1648_));
 sg13g2_or2_1 _4794_ (.X(_1651_),
    .B(_1650_),
    .A(_1644_));
 sg13g2_nand2_1 _4795_ (.Y(_1652_),
    .A(_1644_),
    .B(_1650_));
 sg13g2_and3_1 _4796_ (.X(_0200_),
    .A(net483),
    .B(_1651_),
    .C(_1652_));
 sg13g2_nor3_1 _4797_ (.A(net536),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][12] ),
    .C(_1646_),
    .Y(_1653_));
 sg13g2_o21ai_1 _4798_ (.B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][12] ),
    .Y(_1654_),
    .A1(net536),
    .A2(_1646_));
 sg13g2_nor2b_1 _4799_ (.A(_1653_),
    .B_N(_1654_),
    .Y(_1655_));
 sg13g2_nand2_1 _4800_ (.Y(_1656_),
    .A(net1383),
    .B(_1655_));
 sg13g2_xnor2_1 _4801_ (.Y(_1657_),
    .A(net1383),
    .B(_1655_));
 sg13g2_nand3_1 _4802_ (.B(_1652_),
    .C(_1657_),
    .A(_1649_),
    .Y(_1658_));
 sg13g2_a21o_1 _4803_ (.A2(_1652_),
    .A1(_1649_),
    .B1(_1657_),
    .X(_1659_));
 sg13g2_and3_1 _4804_ (.X(_0201_),
    .A(net483),
    .B(_1658_),
    .C(_1659_));
 sg13g2_a21oi_2 _4805_ (.B1(_1653_),
    .Y(_1660_),
    .A2(net1569),
    .A1(net536));
 sg13g2_nand2_1 _4806_ (.Y(_1661_),
    .A(net1237),
    .B(net391));
 sg13g2_xnor2_1 _4807_ (.Y(_1662_),
    .A(net1237),
    .B(net392));
 sg13g2_nand3_1 _4808_ (.B(_1659_),
    .C(_1662_),
    .A(_1656_),
    .Y(_1663_));
 sg13g2_a21o_2 _4809_ (.A2(_1659_),
    .A1(_1656_),
    .B1(_1662_),
    .X(_1664_));
 sg13g2_and3_1 _4810_ (.X(_0202_),
    .A(net471),
    .B(_1663_),
    .C(_1664_));
 sg13g2_xnor2_1 _4811_ (.Y(_1665_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][5] ),
    .B(net391));
 sg13g2_a21oi_1 _4812_ (.A1(_1661_),
    .A2(_1664_),
    .Y(_1666_),
    .B1(_1665_));
 sg13g2_and3_1 _4813_ (.X(_1667_),
    .A(_1661_),
    .B(_1664_),
    .C(_1665_));
 sg13g2_nor3_1 _4814_ (.A(net426),
    .B(net1238),
    .C(_1667_),
    .Y(_0203_));
 sg13g2_o21ai_1 _4815_ (.B1(net391),
    .Y(_1668_),
    .A1(net1237),
    .A2(net1545));
 sg13g2_o21ai_1 _4816_ (.B1(_1668_),
    .Y(_1669_),
    .A1(_1664_),
    .A2(_1665_));
 sg13g2_xnor2_1 _4817_ (.Y(_1670_),
    .A(net1091),
    .B(net391));
 sg13g2_inv_1 _4818_ (.Y(_1671_),
    .A(_1670_));
 sg13g2_and2_1 _4819_ (.A(_1669_),
    .B(_1671_),
    .X(_1672_));
 sg13g2_o21ai_1 _4820_ (.B1(net468),
    .Y(_1673_),
    .A1(_1669_),
    .A2(_1671_));
 sg13g2_nor2_1 _4821_ (.A(_1672_),
    .B(_1673_),
    .Y(_0204_));
 sg13g2_a21oi_1 _4822_ (.A1(net1091),
    .A2(net391),
    .Y(_1674_),
    .B1(_1672_));
 sg13g2_xnor2_1 _4823_ (.Y(_1675_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][7] ),
    .B(net391));
 sg13g2_o21ai_1 _4824_ (.B1(net468),
    .Y(_1676_),
    .A1(_1674_),
    .A2(_1675_));
 sg13g2_a21oi_1 _4825_ (.A1(_1674_),
    .A2(_1675_),
    .Y(_0205_),
    .B1(_1676_));
 sg13g2_o21ai_1 _4826_ (.B1(_1671_),
    .Y(_1677_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][7] ),
    .A2(net391));
 sg13g2_or3_1 _4827_ (.A(_1664_),
    .B(_1665_),
    .C(_1677_),
    .X(_1678_));
 sg13g2_o21ai_1 _4828_ (.B1(net391),
    .Y(_1679_),
    .A1(net1091),
    .A2(net1515));
 sg13g2_nand3_1 _4829_ (.B(_1678_),
    .C(_1679_),
    .A(_1668_),
    .Y(_1680_));
 sg13g2_xnor2_1 _4830_ (.Y(_1681_),
    .A(net1137),
    .B(net392));
 sg13g2_nor2b_1 _4831_ (.A(net1516),
    .B_N(_1681_),
    .Y(_1682_));
 sg13g2_nor2b_1 _4832_ (.A(_1681_),
    .B_N(_1680_),
    .Y(_1683_));
 sg13g2_nor3_1 _4833_ (.A(net426),
    .B(_1682_),
    .C(_1683_),
    .Y(_0206_));
 sg13g2_xnor2_1 _4834_ (.Y(_1684_),
    .A(net1044),
    .B(_1660_));
 sg13g2_inv_1 _4835_ (.Y(_1685_),
    .A(_1684_));
 sg13g2_a21oi_1 _4836_ (.A1(net1137),
    .A2(net392),
    .Y(_1686_),
    .B1(_1683_));
 sg13g2_o21ai_1 _4837_ (.B1(net471),
    .Y(_1687_),
    .A1(_1684_),
    .A2(_1686_));
 sg13g2_a21oi_1 _4838_ (.A1(_1684_),
    .A2(_1686_),
    .Y(_0207_),
    .B1(_1687_));
 sg13g2_nand2_1 _4839_ (.Y(_1688_),
    .A(net1261),
    .B(_1660_));
 sg13g2_xnor2_1 _4840_ (.Y(_1689_),
    .A(net1261),
    .B(net392));
 sg13g2_nand2_1 _4841_ (.Y(_1690_),
    .A(_1683_),
    .B(_1685_));
 sg13g2_o21ai_1 _4842_ (.B1(net392),
    .Y(_1691_),
    .A1(net1044),
    .A2(net1137));
 sg13g2_nand3_1 _4843_ (.B(_1690_),
    .C(_1691_),
    .A(_1689_),
    .Y(_1692_));
 sg13g2_a21o_1 _4844_ (.A2(_1691_),
    .A1(_1690_),
    .B1(_1689_),
    .X(_1693_));
 sg13g2_and3_1 _4845_ (.X(_0208_),
    .A(net471),
    .B(_1692_),
    .C(_1693_));
 sg13g2_xnor2_1 _4846_ (.Y(_1694_),
    .A(net1201),
    .B(net392));
 sg13g2_and2_1 _4847_ (.A(_1688_),
    .B(_1693_),
    .X(_1695_));
 sg13g2_o21ai_1 _4848_ (.B1(net471),
    .Y(_1696_),
    .A1(_1694_),
    .A2(_1695_));
 sg13g2_a21oi_1 _4849_ (.A1(_1694_),
    .A2(_1695_),
    .Y(_0209_),
    .B1(_1696_));
 sg13g2_or3_1 _4850_ (.A(_1689_),
    .B(_1690_),
    .C(_1694_),
    .X(_1697_));
 sg13g2_o21ai_1 _4851_ (.B1(net392),
    .Y(_1698_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[1] ),
    .A2(net1201));
 sg13g2_nand3_1 _4852_ (.B(_1697_),
    .C(net1202),
    .A(_1691_),
    .Y(_1699_));
 sg13g2_xor2_1 _4853_ (.B(_1660_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[10] ),
    .X(_1700_));
 sg13g2_o21ai_1 _4854_ (.B1(net483),
    .Y(_1701_),
    .A1(_1699_),
    .A2(_1700_));
 sg13g2_a21oi_1 _4855_ (.A1(_1699_),
    .A2(_1700_),
    .Y(_0210_),
    .B1(_1701_));
 sg13g2_nand2_1 _4856_ (.Y(_1702_),
    .A(net998),
    .B(net1044));
 sg13g2_o21ai_1 _4857_ (.B1(net483),
    .Y(_1703_),
    .A1(net998),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[0] ));
 sg13g2_nor2b_1 _4858_ (.A(net999),
    .B_N(_1702_),
    .Y(_0211_));
 sg13g2_nor2b_1 _4859_ (.A(net536),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[0] ),
    .Y(_1704_));
 sg13g2_xnor2_1 _4860_ (.Y(_1705_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[1] ),
    .B(_1704_));
 sg13g2_or2_1 _4861_ (.X(_1706_),
    .B(_1705_),
    .A(_0614_));
 sg13g2_xnor2_1 _4862_ (.Y(_1707_),
    .A(_0614_),
    .B(_1705_));
 sg13g2_o21ai_1 _4863_ (.B1(net483),
    .Y(_1708_),
    .A1(_1702_),
    .A2(_1707_));
 sg13g2_a21oi_1 _4864_ (.A1(_1702_),
    .A2(_1707_),
    .Y(_0212_),
    .B1(_1708_));
 sg13g2_o21ai_1 _4865_ (.B1(_1706_),
    .Y(_1709_),
    .A1(_1702_),
    .A2(_1707_));
 sg13g2_o21ai_1 _4866_ (.B1(_0613_),
    .Y(_1710_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[0] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[1] ));
 sg13g2_xnor2_1 _4867_ (.Y(_1711_),
    .A(_0615_),
    .B(_1710_));
 sg13g2_xnor2_1 _4868_ (.Y(_1712_),
    .A(_0616_),
    .B(_1711_));
 sg13g2_nand2b_1 _4869_ (.Y(_1713_),
    .B(_1712_),
    .A_N(_1709_));
 sg13g2_nand2b_1 _4870_ (.Y(_1714_),
    .B(_1709_),
    .A_N(_1712_));
 sg13g2_and3_1 _4871_ (.X(_0213_),
    .A(net484),
    .B(_1713_),
    .C(_1714_));
 sg13g2_o21ai_1 _4872_ (.B1(_1714_),
    .Y(_1715_),
    .A1(_0616_),
    .A2(_1711_));
 sg13g2_a21oi_1 _4873_ (.A1(_0615_),
    .A2(_1710_),
    .Y(_1716_),
    .B1(net536));
 sg13g2_xnor2_1 _4874_ (.Y(_1717_),
    .A(net1493),
    .B(_1716_));
 sg13g2_nor2b_1 _4875_ (.A(_1717_),
    .B_N(net1447),
    .Y(_1718_));
 sg13g2_xnor2_1 _4876_ (.Y(_1719_),
    .A(net1447),
    .B(_1717_));
 sg13g2_o21ai_1 _4877_ (.B1(net483),
    .Y(_1720_),
    .A1(_1715_),
    .A2(_1719_));
 sg13g2_a21oi_1 _4878_ (.A1(_1715_),
    .A2(_1719_),
    .Y(_0214_),
    .B1(_1720_));
 sg13g2_a21oi_2 _4879_ (.B1(_1718_),
    .Y(_1721_),
    .A2(_1719_),
    .A1(_1715_));
 sg13g2_mux2_1 _4880_ (.A0(_1716_),
    .A1(net536),
    .S(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[10] ),
    .X(_1722_));
 sg13g2_xnor2_1 _4881_ (.Y(_1723_),
    .A(net1167),
    .B(net389));
 sg13g2_nor2_1 _4882_ (.A(_1721_),
    .B(_1723_),
    .Y(_1724_));
 sg13g2_o21ai_1 _4883_ (.B1(net484),
    .Y(_1725_),
    .A1(_1721_),
    .A2(_1723_));
 sg13g2_a21oi_1 _4884_ (.A1(_1721_),
    .A2(_1723_),
    .Y(_0215_),
    .B1(_1725_));
 sg13g2_a21oi_1 _4885_ (.A1(net1167),
    .A2(net389),
    .Y(_1726_),
    .B1(_1724_));
 sg13g2_xor2_1 _4886_ (.B(net389),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][5] ),
    .X(_1727_));
 sg13g2_inv_1 _4887_ (.Y(_1728_),
    .A(_1727_));
 sg13g2_o21ai_1 _4888_ (.B1(net485),
    .Y(_1729_),
    .A1(_1726_),
    .A2(_1728_));
 sg13g2_a21oi_1 _4889_ (.A1(_1726_),
    .A2(_1728_),
    .Y(_0216_),
    .B1(_1729_));
 sg13g2_nand2_1 _4890_ (.Y(_1730_),
    .A(_1724_),
    .B(_1727_));
 sg13g2_o21ai_1 _4891_ (.B1(net389),
    .Y(_1731_),
    .A1(net1167),
    .A2(net1533));
 sg13g2_nand2_1 _4892_ (.Y(_1732_),
    .A(_1730_),
    .B(_1731_));
 sg13g2_nand2_1 _4893_ (.Y(_1733_),
    .A(net1251),
    .B(net389));
 sg13g2_xor2_1 _4894_ (.B(net389),
    .A(net1251),
    .X(_1734_));
 sg13g2_nand2_1 _4895_ (.Y(_1735_),
    .A(_1732_),
    .B(_1734_));
 sg13g2_o21ai_1 _4896_ (.B1(net485),
    .Y(_1736_),
    .A1(_1732_),
    .A2(_1734_));
 sg13g2_nor2b_1 _4897_ (.A(_1736_),
    .B_N(_1735_),
    .Y(_0217_));
 sg13g2_nand2_1 _4898_ (.Y(_1737_),
    .A(_1733_),
    .B(_1735_));
 sg13g2_xor2_1 _4899_ (.B(net390),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][7] ),
    .X(_1738_));
 sg13g2_o21ai_1 _4900_ (.B1(net485),
    .Y(_1739_),
    .A1(_1737_),
    .A2(_1738_));
 sg13g2_a21oi_1 _4901_ (.A1(_1737_),
    .A2(_1738_),
    .Y(_0218_),
    .B1(_1739_));
 sg13g2_o21ai_1 _4902_ (.B1(_1734_),
    .Y(_1740_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][7] ),
    .A2(net389));
 sg13g2_nor4_1 _4903_ (.A(_1721_),
    .B(_1723_),
    .C(_1728_),
    .D(_1740_),
    .Y(_1741_));
 sg13g2_o21ai_1 _4904_ (.B1(net389),
    .Y(_1742_),
    .A1(net1432),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][7] ));
 sg13g2_nand2_1 _4905_ (.Y(_1743_),
    .A(_1731_),
    .B(_1742_));
 sg13g2_nor2_1 _4906_ (.A(_1741_),
    .B(_1743_),
    .Y(_1744_));
 sg13g2_nand2_1 _4907_ (.Y(_1745_),
    .A(net1173),
    .B(net388));
 sg13g2_xnor2_1 _4908_ (.Y(_1746_),
    .A(net1173),
    .B(net388));
 sg13g2_or2_1 _4909_ (.X(_1747_),
    .B(_1746_),
    .A(_1744_));
 sg13g2_nand2_1 _4910_ (.Y(_1748_),
    .A(net484),
    .B(_1747_));
 sg13g2_a21oi_1 _4911_ (.A1(_1744_),
    .A2(_1746_),
    .Y(_0219_),
    .B1(_1748_));
 sg13g2_xor2_1 _4912_ (.B(net390),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][9] ),
    .X(_1749_));
 sg13g2_nand2_1 _4913_ (.Y(_1750_),
    .A(_1745_),
    .B(_1747_));
 sg13g2_o21ai_1 _4914_ (.B1(net484),
    .Y(_1751_),
    .A1(_1749_),
    .A2(_1750_));
 sg13g2_a21oi_1 _4915_ (.A1(_1749_),
    .A2(_1750_),
    .Y(_0220_),
    .B1(_1751_));
 sg13g2_nand2_1 _4916_ (.Y(_1752_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][10] ),
    .B(net388));
 sg13g2_xor2_1 _4917_ (.B(net388),
    .A(net1564),
    .X(_1753_));
 sg13g2_nor2b_1 _4918_ (.A(_1747_),
    .B_N(_1749_),
    .Y(_1754_));
 sg13g2_o21ai_1 _4919_ (.B1(net388),
    .Y(_1755_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][9] ),
    .A2(net1173));
 sg13g2_inv_1 _4920_ (.Y(_1756_),
    .A(_1755_));
 sg13g2_nor3_1 _4921_ (.A(_1753_),
    .B(_1754_),
    .C(_1756_),
    .Y(_1757_));
 sg13g2_o21ai_1 _4922_ (.B1(_1753_),
    .Y(_1758_),
    .A1(_1754_),
    .A2(_1756_));
 sg13g2_nand2_1 _4923_ (.Y(_1759_),
    .A(net483),
    .B(_1758_));
 sg13g2_nor2_1 _4924_ (.A(net1565),
    .B(_1759_),
    .Y(_0221_));
 sg13g2_xor2_1 _4925_ (.B(net388),
    .A(net1341),
    .X(_1760_));
 sg13g2_inv_1 _4926_ (.Y(_1761_),
    .A(_1760_));
 sg13g2_and2_1 _4927_ (.A(_1752_),
    .B(_1758_),
    .X(_1762_));
 sg13g2_o21ai_1 _4928_ (.B1(net484),
    .Y(_1763_),
    .A1(_1761_),
    .A2(_1762_));
 sg13g2_a21oi_1 _4929_ (.A1(_1761_),
    .A2(_1762_),
    .Y(_0222_),
    .B1(_1763_));
 sg13g2_nand3_1 _4930_ (.B(_1754_),
    .C(_1760_),
    .A(_1753_),
    .Y(_1764_));
 sg13g2_o21ai_1 _4931_ (.B1(net388),
    .Y(_1765_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][10] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][11] ));
 sg13g2_and3_1 _4932_ (.X(_1766_),
    .A(_1755_),
    .B(_1764_),
    .C(_1765_));
 sg13g2_xnor2_1 _4933_ (.Y(_1767_),
    .A(net1215),
    .B(net388));
 sg13g2_o21ai_1 _4934_ (.B1(net483),
    .Y(_1768_),
    .A1(_1766_),
    .A2(_1767_));
 sg13g2_a21oi_1 _4935_ (.A1(_1766_),
    .A2(_1767_),
    .Y(_0223_),
    .B1(_1768_));
 sg13g2_nor2_1 _4936_ (.A(net946),
    .B(_0544_),
    .Y(_1769_));
 sg13g2_xnor2_1 _4937_ (.Y(_1770_),
    .A(net946),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][10] ));
 sg13g2_nor2_1 _4938_ (.A(net426),
    .B(net947),
    .Y(_0224_));
 sg13g2_nor2b_1 _4939_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].z_sign ),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][10] ),
    .Y(_1771_));
 sg13g2_xnor2_1 _4940_ (.Y(_1772_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][11] ),
    .B(_1771_));
 sg13g2_nand2_1 _4941_ (.Y(_1773_),
    .A(net1160),
    .B(_1772_));
 sg13g2_xnor2_1 _4942_ (.Y(_1774_),
    .A(net1160),
    .B(_1772_));
 sg13g2_o21ai_1 _4943_ (.B1(net469),
    .Y(_1775_),
    .A1(_1769_),
    .A2(_1774_));
 sg13g2_a21oi_1 _4944_ (.A1(_1769_),
    .A2(_1774_),
    .Y(_0225_),
    .B1(_1775_));
 sg13g2_o21ai_1 _4945_ (.B1(_1773_),
    .Y(_1776_),
    .A1(_1769_),
    .A2(_1774_));
 sg13g2_o21ai_1 _4946_ (.B1(_0617_),
    .Y(_1777_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][10] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][11] ));
 sg13g2_xor2_1 _4947_ (.B(_1777_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][12] ),
    .X(_1778_));
 sg13g2_nand2_1 _4948_ (.Y(_1779_),
    .A(net1464),
    .B(_1778_));
 sg13g2_xnor2_1 _4949_ (.Y(_1780_),
    .A(net1464),
    .B(_1778_));
 sg13g2_nand2b_1 _4950_ (.Y(_1781_),
    .B(_1780_),
    .A_N(_1776_));
 sg13g2_nand2b_1 _4951_ (.Y(_1782_),
    .B(_1776_),
    .A_N(_1780_));
 sg13g2_and3_1 _4952_ (.X(_0226_),
    .A(net469),
    .B(_1781_),
    .C(_1782_));
 sg13g2_mux2_1 _4953_ (.A0(_1777_),
    .A1(_0617_),
    .S(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][12] ),
    .X(_1783_));
 sg13g2_or2_1 _4954_ (.X(_1784_),
    .B(net399),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][3] ));
 sg13g2_xnor2_1 _4955_ (.Y(_1785_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][3] ),
    .B(net399));
 sg13g2_nand3_1 _4956_ (.B(_1782_),
    .C(_1785_),
    .A(_1779_),
    .Y(_1786_));
 sg13g2_a21o_1 _4957_ (.A2(_1782_),
    .A1(_1779_),
    .B1(_1785_),
    .X(_1787_));
 sg13g2_and3_1 _4958_ (.X(_0227_),
    .A(net464),
    .B(net1465),
    .C(_1787_));
 sg13g2_nand3b_1 _4959_ (.B(_1784_),
    .C(_1776_),
    .Y(_1788_),
    .A_N(_1780_));
 sg13g2_a22oi_1 _4960_ (.Y(_1789_),
    .B1(net399),
    .B2(net1494),
    .A2(_1778_),
    .A1(net1464));
 sg13g2_xnor2_1 _4961_ (.Y(_1790_),
    .A(net1112),
    .B(net399));
 sg13g2_nand3_1 _4962_ (.B(_1789_),
    .C(_1790_),
    .A(_1788_),
    .Y(_1791_));
 sg13g2_a21oi_1 _4963_ (.A1(_1788_),
    .A2(_1789_),
    .Y(_1792_),
    .B1(_1790_));
 sg13g2_and2_1 _4964_ (.A(net469),
    .B(_1791_),
    .X(_1793_));
 sg13g2_nor2b_1 _4965_ (.A(_1792_),
    .B_N(_1793_),
    .Y(_0228_));
 sg13g2_a21oi_1 _4966_ (.A1(net1112),
    .A2(net398),
    .Y(_1794_),
    .B1(_1792_));
 sg13g2_xnor2_1 _4967_ (.Y(_1795_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][5] ),
    .B(net397));
 sg13g2_inv_1 _4968_ (.Y(_1796_),
    .A(_1795_));
 sg13g2_o21ai_1 _4969_ (.B1(net467),
    .Y(_1797_),
    .A1(_1794_),
    .A2(_1795_));
 sg13g2_a21oi_1 _4970_ (.A1(_1794_),
    .A2(_1795_),
    .Y(_0229_),
    .B1(_1797_));
 sg13g2_nand2_1 _4971_ (.Y(_1798_),
    .A(_1792_),
    .B(_1796_));
 sg13g2_o21ai_1 _4972_ (.B1(net397),
    .Y(_1799_),
    .A1(net1543),
    .A2(net1573));
 sg13g2_and2_1 _4973_ (.A(_1798_),
    .B(net1544),
    .X(_1800_));
 sg13g2_xnor2_1 _4974_ (.Y(_1801_),
    .A(net1122),
    .B(net397));
 sg13g2_nor2_1 _4975_ (.A(_1800_),
    .B(_1801_),
    .Y(_1802_));
 sg13g2_a21oi_1 _4976_ (.A1(_1800_),
    .A2(_1801_),
    .Y(_1803_),
    .B1(net426));
 sg13g2_nor2b_1 _4977_ (.A(_1802_),
    .B_N(_1803_),
    .Y(_0230_));
 sg13g2_a21oi_1 _4978_ (.A1(net1122),
    .A2(net397),
    .Y(_1804_),
    .B1(_1802_));
 sg13g2_xnor2_1 _4979_ (.Y(_1805_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][7] ),
    .B(net397));
 sg13g2_o21ai_1 _4980_ (.B1(net467),
    .Y(_1806_),
    .A1(_1804_),
    .A2(_1805_));
 sg13g2_a21oi_1 _4981_ (.A1(_1804_),
    .A2(_1805_),
    .Y(_0231_),
    .B1(_1806_));
 sg13g2_nor2_1 _4982_ (.A(_1798_),
    .B(_1801_),
    .Y(_1807_));
 sg13g2_o21ai_1 _4983_ (.B1(_1807_),
    .Y(_1808_),
    .A1(net1433),
    .A2(net397));
 sg13g2_o21ai_1 _4984_ (.B1(net397),
    .Y(_1809_),
    .A1(net1122),
    .A2(net1433));
 sg13g2_and3_1 _4985_ (.X(_1810_),
    .A(_1799_),
    .B(_1808_),
    .C(_1809_));
 sg13g2_nand2_1 _4986_ (.Y(_1811_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][8] ),
    .B(net397));
 sg13g2_xnor2_1 _4987_ (.Y(_1812_),
    .A(net1421),
    .B(net398));
 sg13g2_o21ai_1 _4988_ (.B1(net468),
    .Y(_1813_),
    .A1(_1810_),
    .A2(_1812_));
 sg13g2_a21oi_1 _4989_ (.A1(net1434),
    .A2(_1812_),
    .Y(_0232_),
    .B1(_1813_));
 sg13g2_o21ai_1 _4990_ (.B1(_1811_),
    .Y(_1814_),
    .A1(_1810_),
    .A2(_1812_));
 sg13g2_nand2_1 _4991_ (.Y(_1815_),
    .A(net1186),
    .B(net398));
 sg13g2_xor2_1 _4992_ (.B(net398),
    .A(net1186),
    .X(_1816_));
 sg13g2_o21ai_1 _4993_ (.B1(net468),
    .Y(_1817_),
    .A1(_1814_),
    .A2(_1816_));
 sg13g2_a21oi_1 _4994_ (.A1(_1814_),
    .A2(_1816_),
    .Y(_0233_),
    .B1(_1817_));
 sg13g2_xnor2_1 _4995_ (.Y(_1818_),
    .A(net1052),
    .B(net399));
 sg13g2_o21ai_1 _4996_ (.B1(_1814_),
    .Y(_1819_),
    .A1(net1186),
    .A2(net398));
 sg13g2_and3_1 _4997_ (.X(_1820_),
    .A(_1815_),
    .B(_1818_),
    .C(_1819_));
 sg13g2_a21oi_1 _4998_ (.A1(_1815_),
    .A2(_1819_),
    .Y(_1821_),
    .B1(_1818_));
 sg13g2_nor3_1 _4999_ (.A(net426),
    .B(_1820_),
    .C(_1821_),
    .Y(_0234_));
 sg13g2_a21oi_1 _5000_ (.A1(net1052),
    .A2(net399),
    .Y(_1822_),
    .B1(_1821_));
 sg13g2_xnor2_1 _5001_ (.Y(_1823_),
    .A(net1196),
    .B(net399));
 sg13g2_o21ai_1 _5002_ (.B1(net469),
    .Y(_1824_),
    .A1(_1822_),
    .A2(_1823_));
 sg13g2_a21oi_1 _5003_ (.A1(_1822_),
    .A2(_1823_),
    .Y(_0235_),
    .B1(_1824_));
 sg13g2_nand2_1 _5004_ (.Y(_1825_),
    .A(net988),
    .B(net1052));
 sg13g2_o21ai_1 _5005_ (.B1(net469),
    .Y(_1826_),
    .A1(net988),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[0] ));
 sg13g2_nor2b_1 _5006_ (.A(net989),
    .B_N(_1825_),
    .Y(_0236_));
 sg13g2_nand2_1 _5007_ (.Y(_1827_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[0] ),
    .B(_0617_));
 sg13g2_xnor2_1 _5008_ (.Y(_1828_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[1] ),
    .B(_1827_));
 sg13g2_nand2_1 _5009_ (.Y(_1829_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][1] ),
    .B(_1828_));
 sg13g2_xnor2_1 _5010_ (.Y(_1830_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][1] ),
    .B(_1828_));
 sg13g2_o21ai_1 _5011_ (.B1(net469),
    .Y(_1831_),
    .A1(_1825_),
    .A2(_1830_));
 sg13g2_a21oi_1 _5012_ (.A1(_1825_),
    .A2(_1830_),
    .Y(_0237_),
    .B1(_1831_));
 sg13g2_o21ai_1 _5013_ (.B1(_1829_),
    .Y(_1832_),
    .A1(_1825_),
    .A2(_1830_));
 sg13g2_nor2_1 _5014_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[0] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[1] ),
    .Y(_1833_));
 sg13g2_nor3_1 _5015_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].z_sign ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[10] ),
    .C(_1833_),
    .Y(_1834_));
 sg13g2_o21ai_1 _5016_ (.B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[10] ),
    .Y(_1835_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].z_sign ),
    .A2(_1833_));
 sg13g2_nor2b_1 _5017_ (.A(_1834_),
    .B_N(_1835_),
    .Y(_1836_));
 sg13g2_nor2b_1 _5018_ (.A(_1836_),
    .B_N(net1488),
    .Y(_1837_));
 sg13g2_xnor2_1 _5019_ (.Y(_1838_),
    .A(net1488),
    .B(_1836_));
 sg13g2_nor2_1 _5020_ (.A(_1832_),
    .B(_1838_),
    .Y(_1839_));
 sg13g2_a21oi_1 _5021_ (.A1(_1832_),
    .A2(_1838_),
    .Y(_1840_),
    .B1(net427));
 sg13g2_nor2b_1 _5022_ (.A(net1489),
    .B_N(_1840_),
    .Y(_0238_));
 sg13g2_a21oi_1 _5023_ (.A1(_1832_),
    .A2(_1838_),
    .Y(_1841_),
    .B1(_1837_));
 sg13g2_a21oi_2 _5024_ (.B1(_1834_),
    .Y(_1842_),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[10] ),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].z_sign ));
 sg13g2_a21o_2 _5025_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[10] ),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].z_sign ),
    .B1(_1834_),
    .X(_1843_));
 sg13g2_nand2_1 _5026_ (.Y(_1844_),
    .A(net1500),
    .B(net395));
 sg13g2_xnor2_1 _5027_ (.Y(_1845_),
    .A(net1500),
    .B(net396));
 sg13g2_nand2b_1 _5028_ (.Y(_1846_),
    .B(_1841_),
    .A_N(_1845_));
 sg13g2_nand2b_1 _5029_ (.Y(_1847_),
    .B(_1845_),
    .A_N(_1841_));
 sg13g2_and3_1 _5030_ (.X(_0239_),
    .A(net470),
    .B(_1846_),
    .C(_1847_));
 sg13g2_xnor2_1 _5031_ (.Y(_1848_),
    .A(_0618_),
    .B(_1842_));
 sg13g2_nand3_1 _5032_ (.B(_1847_),
    .C(_1848_),
    .A(_1844_),
    .Y(_1849_));
 sg13g2_a21o_2 _5033_ (.A2(_1847_),
    .A1(_1844_),
    .B1(_1848_),
    .X(_1850_));
 sg13g2_and3_1 _5034_ (.X(_0240_),
    .A(net470),
    .B(_1849_),
    .C(_1850_));
 sg13g2_o21ai_1 _5035_ (.B1(_1850_),
    .Y(_1851_),
    .A1(_0618_),
    .A2(net396));
 sg13g2_xnor2_1 _5036_ (.Y(_1852_),
    .A(net1396),
    .B(net396));
 sg13g2_inv_1 _5037_ (.Y(_1853_),
    .A(_1852_));
 sg13g2_o21ai_1 _5038_ (.B1(net470),
    .Y(_1854_),
    .A1(_1851_),
    .A2(_1852_));
 sg13g2_a21oi_1 _5039_ (.A1(_1851_),
    .A2(_1852_),
    .Y(_0241_),
    .B1(_1854_));
 sg13g2_o21ai_1 _5040_ (.B1(net395),
    .Y(_1855_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][4] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][5] ));
 sg13g2_o21ai_1 _5041_ (.B1(_1855_),
    .Y(_1856_),
    .A1(_1850_),
    .A2(_1853_));
 sg13g2_nand2_1 _5042_ (.Y(_1857_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][6] ),
    .B(_1843_));
 sg13g2_xnor2_1 _5043_ (.Y(_1858_),
    .A(net1560),
    .B(net396));
 sg13g2_nand2_1 _5044_ (.Y(_1859_),
    .A(_1856_),
    .B(_1858_));
 sg13g2_o21ai_1 _5045_ (.B1(net470),
    .Y(_1860_),
    .A1(_1856_),
    .A2(_1858_));
 sg13g2_nor2b_2 _5046_ (.A(_1860_),
    .B_N(_1859_),
    .Y(_0242_));
 sg13g2_nand2_1 _5047_ (.Y(_1861_),
    .A(_1857_),
    .B(_1859_));
 sg13g2_xnor2_1 _5048_ (.Y(_1862_),
    .A(net1430),
    .B(net396));
 sg13g2_o21ai_1 _5049_ (.B1(net464),
    .Y(_1863_),
    .A1(_1861_),
    .A2(_1862_));
 sg13g2_a21oi_1 _5050_ (.A1(_1861_),
    .A2(_1862_),
    .Y(_0243_),
    .B1(_1863_));
 sg13g2_o21ai_1 _5051_ (.B1(_1858_),
    .Y(_1864_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][7] ),
    .A2(net395));
 sg13g2_or3_1 _5052_ (.A(_1850_),
    .B(_1853_),
    .C(_1864_),
    .X(_1865_));
 sg13g2_nand2_1 _5053_ (.Y(_1866_),
    .A(_1855_),
    .B(_1857_));
 sg13g2_a21oi_1 _5054_ (.A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][7] ),
    .A2(_1843_),
    .Y(_1867_),
    .B1(_1866_));
 sg13g2_xnor2_1 _5055_ (.Y(_1868_),
    .A(net1219),
    .B(net395));
 sg13g2_and3_1 _5056_ (.X(_1869_),
    .A(_1865_),
    .B(_1867_),
    .C(_1868_));
 sg13g2_a21oi_1 _5057_ (.A1(_1865_),
    .A2(_1867_),
    .Y(_1870_),
    .B1(_1868_));
 sg13g2_nor3_1 _5058_ (.A(net426),
    .B(_1869_),
    .C(net1220),
    .Y(_0244_));
 sg13g2_a21oi_1 _5059_ (.A1(net1219),
    .A2(net395),
    .Y(_1871_),
    .B1(_1870_));
 sg13g2_nand2_1 _5060_ (.Y(_1872_),
    .A(net1260),
    .B(net395));
 sg13g2_nor2_1 _5061_ (.A(net1260),
    .B(net395),
    .Y(_1873_));
 sg13g2_xnor2_1 _5062_ (.Y(_1874_),
    .A(net1260),
    .B(net395));
 sg13g2_o21ai_1 _5063_ (.B1(net465),
    .Y(_1875_),
    .A1(_1871_),
    .A2(_1874_));
 sg13g2_a21oi_1 _5064_ (.A1(_1871_),
    .A2(_1874_),
    .Y(_0245_),
    .B1(_1875_));
 sg13g2_xnor2_1 _5065_ (.Y(_1876_),
    .A(net1548),
    .B(net396));
 sg13g2_o21ai_1 _5066_ (.B1(_1872_),
    .Y(_1877_),
    .A1(_1871_),
    .A2(_1873_));
 sg13g2_nand2_1 _5067_ (.Y(_1878_),
    .A(_1876_),
    .B(_1877_));
 sg13g2_o21ai_1 _5068_ (.B1(net464),
    .Y(_1879_),
    .A1(_1876_),
    .A2(_1877_));
 sg13g2_nor2b_1 _5069_ (.A(_1879_),
    .B_N(_1878_),
    .Y(_0246_));
 sg13g2_o21ai_1 _5070_ (.B1(_1878_),
    .Y(_1880_),
    .A1(_0544_),
    .A2(net396));
 sg13g2_xnor2_1 _5071_ (.Y(_1881_),
    .A(net1197),
    .B(net396));
 sg13g2_o21ai_1 _5072_ (.B1(net464),
    .Y(_1882_),
    .A1(_1880_),
    .A2(_1881_));
 sg13g2_a21oi_1 _5073_ (.A1(_1880_),
    .A2(_1881_),
    .Y(_0247_),
    .B1(_1882_));
 sg13g2_and2_1 _5074_ (.A(net448),
    .B(net2),
    .X(_0248_));
 sg13g2_and2_1 _5075_ (.A(net448),
    .B(net3),
    .X(_0249_));
 sg13g2_and2_1 _5076_ (.A(net448),
    .B(net4),
    .X(_0250_));
 sg13g2_and2_1 _5077_ (.A(net448),
    .B(net5),
    .X(_0251_));
 sg13g2_and2_1 _5078_ (.A(net448),
    .B(net6),
    .X(_0252_));
 sg13g2_and2_1 _5079_ (.A(net448),
    .B(net7),
    .X(_0253_));
 sg13g2_and2_1 _5080_ (.A(net448),
    .B(net8),
    .X(_0254_));
 sg13g2_and2_1 _5081_ (.A(net449),
    .B(net9),
    .X(_0255_));
 sg13g2_and2_1 _5082_ (.A(net449),
    .B(net10),
    .X(_0256_));
 sg13g2_and2_1 _5083_ (.A(net449),
    .B(net11),
    .X(_0257_));
 sg13g2_and2_1 _5084_ (.A(net449),
    .B(net12),
    .X(_0258_));
 sg13g2_and2_1 _5085_ (.A(net450),
    .B(net13),
    .X(_0259_));
 sg13g2_and2_1 _5086_ (.A(net450),
    .B(net14),
    .X(_0260_));
 sg13g2_nor2_1 _5087_ (.A(net803),
    .B(net423),
    .Y(_0261_));
 sg13g2_nand2_1 _5088_ (.Y(_1883_),
    .A(net1033),
    .B(net1101));
 sg13g2_o21ai_1 _5089_ (.B1(net478),
    .Y(_1884_),
    .A1(net1033),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[0] ));
 sg13g2_nor2b_1 _5090_ (.A(net1034),
    .B_N(_1883_),
    .Y(_0262_));
 sg13g2_nand2b_1 _5091_ (.Y(_1885_),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[0] ),
    .A_N(net526));
 sg13g2_xnor2_1 _5092_ (.Y(_1886_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[1] ),
    .B(_1885_));
 sg13g2_nand2_1 _5093_ (.Y(_1887_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][1] ),
    .B(_1886_));
 sg13g2_xnor2_1 _5094_ (.Y(_1888_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][1] ),
    .B(_1886_));
 sg13g2_o21ai_1 _5095_ (.B1(net480),
    .Y(_1889_),
    .A1(_1883_),
    .A2(_1888_));
 sg13g2_a21oi_1 _5096_ (.A1(_1883_),
    .A2(_1888_),
    .Y(_0263_),
    .B1(_1889_));
 sg13g2_o21ai_1 _5097_ (.B1(_1887_),
    .Y(_1890_),
    .A1(_1883_),
    .A2(_1888_));
 sg13g2_or2_1 _5098_ (.X(_1891_),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[1] ),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[0] ));
 sg13g2_a21oi_1 _5099_ (.A1(net415),
    .A2(_1891_),
    .Y(_1892_),
    .B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[2] ));
 sg13g2_nand3_1 _5100_ (.B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[2] ),
    .C(_1891_),
    .A(net415),
    .Y(_1893_));
 sg13g2_nor2b_1 _5101_ (.A(_1892_),
    .B_N(_1893_),
    .Y(_1894_));
 sg13g2_and2_1 _5102_ (.A(net1393),
    .B(_1894_),
    .X(_1895_));
 sg13g2_xor2_1 _5103_ (.B(_1894_),
    .A(net1393),
    .X(_1896_));
 sg13g2_nor2_1 _5104_ (.A(_1890_),
    .B(_1896_),
    .Y(_1897_));
 sg13g2_a21oi_1 _5105_ (.A1(_1890_),
    .A2(_1896_),
    .Y(_1898_),
    .B1(net430));
 sg13g2_nor2b_1 _5106_ (.A(net1394),
    .B_N(_1898_),
    .Y(_0264_));
 sg13g2_a21oi_1 _5107_ (.A1(_1890_),
    .A2(_1896_),
    .Y(_1899_),
    .B1(_1895_));
 sg13g2_nor2_1 _5108_ (.A(net526),
    .B(_1892_),
    .Y(_1900_));
 sg13g2_xnor2_1 _5109_ (.Y(_1901_),
    .A(_0565_),
    .B(_1900_));
 sg13g2_nand2_1 _5110_ (.Y(_1902_),
    .A(net1485),
    .B(_1901_));
 sg13g2_xnor2_1 _5111_ (.Y(_1903_),
    .A(net1485),
    .B(_1901_));
 sg13g2_nor2_1 _5112_ (.A(_1899_),
    .B(_1903_),
    .Y(_1904_));
 sg13g2_a21oi_1 _5113_ (.A1(_1899_),
    .A2(_1903_),
    .Y(_1905_),
    .B1(net430));
 sg13g2_nor2b_1 _5114_ (.A(_1904_),
    .B_N(_1905_),
    .Y(_0265_));
 sg13g2_o21ai_1 _5115_ (.B1(_1902_),
    .Y(_1906_),
    .A1(_1899_),
    .A2(_1903_));
 sg13g2_a21oi_1 _5116_ (.A1(_0565_),
    .A2(_1892_),
    .Y(_1907_),
    .B1(net526));
 sg13g2_nor2_1 _5117_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[4] ),
    .B(_1907_),
    .Y(_1908_));
 sg13g2_xor2_1 _5118_ (.B(_1907_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[4] ),
    .X(_1909_));
 sg13g2_nand2_1 _5119_ (.Y(_1910_),
    .A(net1275),
    .B(_1909_));
 sg13g2_inv_1 _5120_ (.Y(_1911_),
    .A(_1910_));
 sg13g2_xnor2_1 _5121_ (.Y(_1912_),
    .A(net1275),
    .B(_1909_));
 sg13g2_inv_1 _5122_ (.Y(_1913_),
    .A(_1912_));
 sg13g2_nand2b_1 _5123_ (.Y(_1914_),
    .B(_1912_),
    .A_N(_1906_));
 sg13g2_nand2_1 _5124_ (.Y(_1915_),
    .A(_1906_),
    .B(_1913_));
 sg13g2_and3_1 _5125_ (.X(_0266_),
    .A(net492),
    .B(_1914_),
    .C(_1915_));
 sg13g2_nand2_1 _5126_ (.Y(_1916_),
    .A(_1910_),
    .B(_1915_));
 sg13g2_nor2_1 _5127_ (.A(net526),
    .B(_1908_),
    .Y(_1917_));
 sg13g2_xnor2_1 _5128_ (.Y(_1918_),
    .A(_0566_),
    .B(_1917_));
 sg13g2_nor2_1 _5129_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][5] ),
    .B(_1918_),
    .Y(_1919_));
 sg13g2_xnor2_1 _5130_ (.Y(_1920_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][5] ),
    .B(_1918_));
 sg13g2_inv_1 _5131_ (.Y(_1921_),
    .A(_1920_));
 sg13g2_o21ai_1 _5132_ (.B1(net492),
    .Y(_1922_),
    .A1(_1916_),
    .A2(_1921_));
 sg13g2_a21oi_1 _5133_ (.A1(_1916_),
    .A2(_1921_),
    .Y(_0267_),
    .B1(_1922_));
 sg13g2_a21oi_1 _5134_ (.A1(_0566_),
    .A2(_1908_),
    .Y(_1923_),
    .B1(net526));
 sg13g2_or2_1 _5135_ (.X(_1924_),
    .B(_1923_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[6] ));
 sg13g2_xor2_1 _5136_ (.B(_1923_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[6] ),
    .X(_1925_));
 sg13g2_xnor2_1 _5137_ (.Y(_1926_),
    .A(net1162),
    .B(_1925_));
 sg13g2_a221oi_1 _5138_ (.B2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][5] ),
    .C1(_1911_),
    .B1(_1918_),
    .A1(_1906_),
    .Y(_1927_),
    .A2(_1913_));
 sg13g2_or2_1 _5139_ (.X(_1928_),
    .B(_1927_),
    .A(_1919_));
 sg13g2_nor2_1 _5140_ (.A(_1926_),
    .B(_1928_),
    .Y(_1929_));
 sg13g2_nand2b_1 _5141_ (.Y(_1930_),
    .B(net493),
    .A_N(_1929_));
 sg13g2_a21oi_1 _5142_ (.A1(net1163),
    .A2(_1928_),
    .Y(_0268_),
    .B1(_1930_));
 sg13g2_a21o_1 _5143_ (.A2(_1925_),
    .A1(net1162),
    .B1(_1929_),
    .X(_1931_));
 sg13g2_nor2_1 _5144_ (.A(net415),
    .B(_0567_),
    .Y(_1932_));
 sg13g2_nor2_1 _5145_ (.A(net527),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[10] ),
    .Y(_1933_));
 sg13g2_a21oi_2 _5146_ (.B1(_1932_),
    .Y(_1934_),
    .A2(_1933_),
    .A1(_1924_));
 sg13g2_inv_1 _5147_ (.Y(_1935_),
    .A(net380));
 sg13g2_o21ai_1 _5148_ (.B1(net380),
    .Y(_1936_),
    .A1(_0567_),
    .A2(_1924_));
 sg13g2_and2_1 _5149_ (.A(net1410),
    .B(_1936_),
    .X(_1937_));
 sg13g2_xnor2_1 _5150_ (.Y(_1938_),
    .A(_0568_),
    .B(_1936_));
 sg13g2_o21ai_1 _5151_ (.B1(net493),
    .Y(_1939_),
    .A1(_1931_),
    .A2(_1938_));
 sg13g2_a21oi_1 _5152_ (.A1(_1931_),
    .A2(_1938_),
    .Y(_0269_),
    .B1(_1939_));
 sg13g2_a21o_1 _5153_ (.A2(_1938_),
    .A1(_1931_),
    .B1(_1937_),
    .X(_1940_));
 sg13g2_xnor2_1 _5154_ (.Y(_1941_),
    .A(net1558),
    .B(net380));
 sg13g2_nand2_1 _5155_ (.Y(_1942_),
    .A(_1940_),
    .B(_1941_));
 sg13g2_o21ai_1 _5156_ (.B1(net493),
    .Y(_1943_),
    .A1(_1940_),
    .A2(_1941_));
 sg13g2_nor2b_1 _5157_ (.A(_1943_),
    .B_N(_1942_),
    .Y(_0270_));
 sg13g2_xnor2_1 _5158_ (.Y(_1944_),
    .A(net1289),
    .B(_1934_));
 sg13g2_o21ai_1 _5159_ (.B1(_1942_),
    .Y(_1945_),
    .A1(_0569_),
    .A2(net380));
 sg13g2_o21ai_1 _5160_ (.B1(net492),
    .Y(_1946_),
    .A1(_1944_),
    .A2(_1945_));
 sg13g2_a21oi_1 _5161_ (.A1(_1944_),
    .A2(_1945_),
    .Y(_0271_),
    .B1(_1946_));
 sg13g2_xnor2_1 _5162_ (.Y(_1947_),
    .A(_0571_),
    .B(net380));
 sg13g2_nand3_1 _5163_ (.B(_1941_),
    .C(_1944_),
    .A(_1940_),
    .Y(_1948_));
 sg13g2_o21ai_1 _5164_ (.B1(_1935_),
    .Y(_1949_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][8] ),
    .A2(net1289));
 sg13g2_nand3_1 _5165_ (.B(_1948_),
    .C(_1949_),
    .A(_1947_),
    .Y(_1950_));
 sg13g2_a21o_1 _5166_ (.A2(_1949_),
    .A1(_1948_),
    .B1(_1947_),
    .X(_1951_));
 sg13g2_and3_1 _5167_ (.X(_0272_),
    .A(net493),
    .B(_1950_),
    .C(_1951_));
 sg13g2_xnor2_1 _5168_ (.Y(_1952_),
    .A(net1291),
    .B(net380));
 sg13g2_o21ai_1 _5169_ (.B1(_1951_),
    .Y(_1953_),
    .A1(_0571_),
    .A2(net380));
 sg13g2_o21ai_1 _5170_ (.B1(net493),
    .Y(_1954_),
    .A1(_1952_),
    .A2(_1953_));
 sg13g2_a21oi_1 _5171_ (.A1(_1952_),
    .A2(_1953_),
    .Y(_0273_),
    .B1(_1954_));
 sg13g2_nor2_1 _5172_ (.A(_1947_),
    .B(_1948_),
    .Y(_1955_));
 sg13g2_o21ai_1 _5173_ (.B1(_1935_),
    .Y(_1956_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][10] ),
    .A2(net1291));
 sg13g2_nand2_1 _5174_ (.Y(_1957_),
    .A(_1949_),
    .B(_1956_));
 sg13g2_a21oi_1 _5175_ (.A1(_1952_),
    .A2(_1955_),
    .Y(_1958_),
    .B1(_1957_));
 sg13g2_xor2_1 _5176_ (.B(net380),
    .A(net1408),
    .X(_1959_));
 sg13g2_o21ai_1 _5177_ (.B1(net492),
    .Y(_1960_),
    .A1(_1958_),
    .A2(_1959_));
 sg13g2_a21oi_1 _5178_ (.A1(_1958_),
    .A2(_1959_),
    .Y(_0274_),
    .B1(_1960_));
 sg13g2_nor2b_1 _5179_ (.A(net912),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][5] ),
    .Y(_1961_));
 sg13g2_xnor2_1 _5180_ (.Y(_1962_),
    .A(net912),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][5] ));
 sg13g2_nor2_1 _5181_ (.A(net439),
    .B(net913),
    .Y(_0275_));
 sg13g2_nor2b_1 _5182_ (.A(net526),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][5] ),
    .Y(_1963_));
 sg13g2_xnor2_1 _5183_ (.Y(_1964_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][6] ),
    .B(_1963_));
 sg13g2_nand2_1 _5184_ (.Y(_1965_),
    .A(net1062),
    .B(_1964_));
 sg13g2_xnor2_1 _5185_ (.Y(_1966_),
    .A(net1062),
    .B(_1964_));
 sg13g2_o21ai_1 _5186_ (.B1(net494),
    .Y(_1967_),
    .A1(_1961_),
    .A2(_1966_));
 sg13g2_a21oi_1 _5187_ (.A1(_1961_),
    .A2(net1063),
    .Y(_0276_),
    .B1(_1967_));
 sg13g2_o21ai_1 _5188_ (.B1(_1965_),
    .Y(_1968_),
    .A1(_1961_),
    .A2(_1966_));
 sg13g2_nor2_1 _5189_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][5] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][6] ),
    .Y(_1969_));
 sg13g2_nor2_1 _5190_ (.A(net527),
    .B(_1969_),
    .Y(_1970_));
 sg13g2_xnor2_1 _5191_ (.Y(_1971_),
    .A(_0568_),
    .B(_1970_));
 sg13g2_nor2b_1 _5192_ (.A(_1971_),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][2] ),
    .Y(_1972_));
 sg13g2_xnor2_1 _5193_ (.Y(_1973_),
    .A(net1337),
    .B(_1971_));
 sg13g2_nor2_1 _5194_ (.A(_1968_),
    .B(_1973_),
    .Y(_1974_));
 sg13g2_a21oi_1 _5195_ (.A1(_1968_),
    .A2(_1973_),
    .Y(_1975_),
    .B1(net439));
 sg13g2_nor2b_1 _5196_ (.A(_1974_),
    .B_N(_1975_),
    .Y(_0277_));
 sg13g2_a21oi_1 _5197_ (.A1(_1968_),
    .A2(_1973_),
    .Y(_1976_),
    .B1(_1972_));
 sg13g2_a21oi_1 _5198_ (.A1(_0568_),
    .A2(_1969_),
    .Y(_1977_),
    .B1(net527));
 sg13g2_xnor2_1 _5199_ (.Y(_1978_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][8] ),
    .B(_1977_));
 sg13g2_nand2_1 _5200_ (.Y(_1979_),
    .A(net1245),
    .B(_1978_));
 sg13g2_xor2_1 _5201_ (.B(_1978_),
    .A(net1245),
    .X(_1980_));
 sg13g2_inv_1 _5202_ (.Y(_1981_),
    .A(_1980_));
 sg13g2_o21ai_1 _5203_ (.B1(net494),
    .Y(_1982_),
    .A1(_1976_),
    .A2(_1981_));
 sg13g2_a21oi_1 _5204_ (.A1(_1976_),
    .A2(_1981_),
    .Y(_0278_),
    .B1(_1982_));
 sg13g2_o21ai_1 _5205_ (.B1(_1979_),
    .Y(_1983_),
    .A1(_1976_),
    .A2(_1981_));
 sg13g2_a21oi_1 _5206_ (.A1(net415),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][8] ),
    .Y(_1984_),
    .B1(_1977_));
 sg13g2_xnor2_1 _5207_ (.Y(_1985_),
    .A(_0570_),
    .B(_1984_));
 sg13g2_and2_1 _5208_ (.A(net1380),
    .B(_1985_),
    .X(_1986_));
 sg13g2_xor2_1 _5209_ (.B(_1985_),
    .A(net1380),
    .X(_1987_));
 sg13g2_nor2_1 _5210_ (.A(_1983_),
    .B(_1987_),
    .Y(_1988_));
 sg13g2_and2_1 _5211_ (.A(_1983_),
    .B(_1987_),
    .X(_1989_));
 sg13g2_nor3_1 _5212_ (.A(net439),
    .B(_1988_),
    .C(_1989_),
    .Y(_0279_));
 sg13g2_nor2_1 _5213_ (.A(_1986_),
    .B(_1989_),
    .Y(_1990_));
 sg13g2_a21oi_1 _5214_ (.A1(_0570_),
    .A2(_1984_),
    .Y(_1991_),
    .B1(net527));
 sg13g2_xnor2_1 _5215_ (.Y(_1992_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][10] ),
    .B(_1991_));
 sg13g2_nor2_1 _5216_ (.A(net1101),
    .B(_1992_),
    .Y(_1993_));
 sg13g2_xnor2_1 _5217_ (.Y(_1994_),
    .A(net1101),
    .B(_1992_));
 sg13g2_xnor2_1 _5218_ (.Y(_1995_),
    .A(_1990_),
    .B(_1994_));
 sg13g2_nor2_1 _5219_ (.A(net439),
    .B(_1995_),
    .Y(_0280_));
 sg13g2_nor2_1 _5220_ (.A(net527),
    .B(_0571_),
    .Y(_1996_));
 sg13g2_nor3_1 _5221_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][11] ),
    .B(_1991_),
    .C(_1996_),
    .Y(_1997_));
 sg13g2_o21ai_1 _5222_ (.B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][11] ),
    .Y(_1998_),
    .A1(_1991_),
    .A2(_1996_));
 sg13g2_nand2b_1 _5223_ (.Y(_1999_),
    .B(_1998_),
    .A_N(_1997_));
 sg13g2_xnor2_1 _5224_ (.Y(_2000_),
    .A(net1538),
    .B(_1999_));
 sg13g2_a221oi_1 _5225_ (.B2(net1542),
    .C1(_1986_),
    .B1(_1992_),
    .A1(_1983_),
    .Y(_2001_),
    .A2(_1987_));
 sg13g2_o21ai_1 _5226_ (.B1(_2000_),
    .Y(_2002_),
    .A1(_1993_),
    .A2(_2001_));
 sg13g2_nor3_1 _5227_ (.A(_1993_),
    .B(_2000_),
    .C(_2001_),
    .Y(_2003_));
 sg13g2_nand2_1 _5228_ (.Y(_2004_),
    .A(net492),
    .B(_2002_));
 sg13g2_nor2_1 _5229_ (.A(_2003_),
    .B(_2004_),
    .Y(_0281_));
 sg13g2_a21o_1 _5230_ (.A2(_1999_),
    .A1(net1538),
    .B1(_2003_),
    .X(_2005_));
 sg13g2_nor3_1 _5231_ (.A(net526),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][12] ),
    .C(_1997_),
    .Y(_2006_));
 sg13g2_a21oi_2 _5232_ (.B1(_2006_),
    .Y(_2007_),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][12] ),
    .A1(net526));
 sg13g2_nand2_1 _5233_ (.Y(_2008_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][12] ),
    .B(_1997_));
 sg13g2_and2_1 _5234_ (.A(net379),
    .B(_2008_),
    .X(_2009_));
 sg13g2_and2_1 _5235_ (.A(net1551),
    .B(_2009_),
    .X(_2010_));
 sg13g2_xnor2_1 _5236_ (.Y(_2011_),
    .A(net1551),
    .B(_2009_));
 sg13g2_nor2b_1 _5237_ (.A(_2005_),
    .B_N(_2011_),
    .Y(_2012_));
 sg13g2_nor2b_1 _5238_ (.A(_2011_),
    .B_N(_2005_),
    .Y(_2013_));
 sg13g2_nor3_1 _5239_ (.A(net430),
    .B(net1539),
    .C(_2013_),
    .Y(_0282_));
 sg13g2_nand2_1 _5240_ (.Y(_2014_),
    .A(net1181),
    .B(net379));
 sg13g2_xnor2_1 _5241_ (.Y(_2015_),
    .A(_0565_),
    .B(net379));
 sg13g2_nor3_1 _5242_ (.A(_2010_),
    .B(_2013_),
    .C(_2015_),
    .Y(_2016_));
 sg13g2_o21ai_1 _5243_ (.B1(_2015_),
    .Y(_2017_),
    .A1(_2010_),
    .A2(_2013_));
 sg13g2_nand2_1 _5244_ (.Y(_2018_),
    .A(net492),
    .B(_2017_));
 sg13g2_nor2_1 _5245_ (.A(_2016_),
    .B(_2018_),
    .Y(_0283_));
 sg13g2_xor2_1 _5246_ (.B(net379),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[4] ),
    .X(_2019_));
 sg13g2_nand2_1 _5247_ (.Y(_2020_),
    .A(_2014_),
    .B(_2017_));
 sg13g2_o21ai_1 _5248_ (.B1(net480),
    .Y(_2021_),
    .A1(_2019_),
    .A2(_2020_));
 sg13g2_a21oi_1 _5249_ (.A1(_2019_),
    .A2(_2020_),
    .Y(_0284_),
    .B1(_2021_));
 sg13g2_nand2_1 _5250_ (.Y(_2022_),
    .A(net1227),
    .B(net379));
 sg13g2_xnor2_1 _5251_ (.Y(_2023_),
    .A(net1227),
    .B(net379));
 sg13g2_nand2b_1 _5252_ (.Y(_2024_),
    .B(_2019_),
    .A_N(_2017_));
 sg13g2_o21ai_1 _5253_ (.B1(_2007_),
    .Y(_2025_),
    .A1(net1181),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[4] ));
 sg13g2_nand3_1 _5254_ (.B(_2024_),
    .C(_2025_),
    .A(_2023_),
    .Y(_2026_));
 sg13g2_a21o_1 _5255_ (.A2(_2025_),
    .A1(_2024_),
    .B1(_2023_),
    .X(_2027_));
 sg13g2_and3_1 _5256_ (.X(_0285_),
    .A(net492),
    .B(_2026_),
    .C(_2027_));
 sg13g2_xnor2_1 _5257_ (.Y(_2028_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[6] ),
    .B(net379));
 sg13g2_and3_1 _5258_ (.X(_2029_),
    .A(_2022_),
    .B(_2027_),
    .C(_2028_));
 sg13g2_a21oi_1 _5259_ (.A1(_2022_),
    .A2(_2027_),
    .Y(_2030_),
    .B1(_2028_));
 sg13g2_nor3_1 _5260_ (.A(net430),
    .B(_2029_),
    .C(net1228),
    .Y(_0286_));
 sg13g2_or3_1 _5261_ (.A(_2023_),
    .B(_2024_),
    .C(_2028_),
    .X(_2031_));
 sg13g2_o21ai_1 _5262_ (.B1(net379),
    .Y(_2032_),
    .A1(net1227),
    .A2(net1314));
 sg13g2_nand3_1 _5263_ (.B(_2031_),
    .C(_2032_),
    .A(_2025_),
    .Y(_2033_));
 sg13g2_xnor2_1 _5264_ (.Y(_2034_),
    .A(_0567_),
    .B(_2007_));
 sg13g2_o21ai_1 _5265_ (.B1(net492),
    .Y(_2035_),
    .A1(_2033_),
    .A2(_2034_));
 sg13g2_a21oi_1 _5266_ (.A1(net1315),
    .A2(_2034_),
    .Y(_0287_),
    .B1(_2035_));
 sg13g2_and2_1 _5267_ (.A(net489),
    .B(net772),
    .X(_0288_));
 sg13g2_and2_1 _5268_ (.A(net489),
    .B(net830),
    .X(_0289_));
 sg13g2_nor2_1 _5269_ (.A(net804),
    .B(net435),
    .Y(_0290_));
 sg13g2_nor2b_1 _5270_ (.A(net528),
    .B_N(net862),
    .Y(_2036_));
 sg13g2_xnor2_1 _5271_ (.Y(_2037_),
    .A(net528),
    .B(net862));
 sg13g2_o21ai_1 _5272_ (.B1(net487),
    .Y(_2038_),
    .A1(net804),
    .A2(_2037_));
 sg13g2_a21oi_1 _5273_ (.A1(net804),
    .A2(_2037_),
    .Y(_0291_),
    .B1(_2038_));
 sg13g2_a21oi_1 _5274_ (.A1(net804),
    .A2(_2037_),
    .Y(_2039_),
    .B1(_2036_));
 sg13g2_nand2_1 _5275_ (.Y(_2040_),
    .A(net528),
    .B(net1095));
 sg13g2_xnor2_1 _5276_ (.Y(_2041_),
    .A(net528),
    .B(net1095));
 sg13g2_or2_1 _5277_ (.X(_2042_),
    .B(_2041_),
    .A(_2039_));
 sg13g2_nand2_1 _5278_ (.Y(_2043_),
    .A(net496),
    .B(_2042_));
 sg13g2_a21oi_1 _5279_ (.A1(_2039_),
    .A2(_2041_),
    .Y(_0292_),
    .B1(_2043_));
 sg13g2_nand2_1 _5280_ (.Y(_2044_),
    .A(net415),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][5] ));
 sg13g2_xor2_1 _5281_ (.B(net1473),
    .A(net528),
    .X(_2045_));
 sg13g2_nand3_1 _5282_ (.B(_2042_),
    .C(_2045_),
    .A(_2040_),
    .Y(_2046_));
 sg13g2_a21o_1 _5283_ (.A2(_2042_),
    .A1(_2040_),
    .B1(_2045_),
    .X(_2047_));
 sg13g2_and3_1 _5284_ (.X(_0293_),
    .A(net496),
    .B(_2046_),
    .C(_2047_));
 sg13g2_and2_1 _5285_ (.A(_2044_),
    .B(_2047_),
    .X(_2048_));
 sg13g2_nand2_1 _5286_ (.Y(_2049_),
    .A(net415),
    .B(net1144));
 sg13g2_xor2_1 _5287_ (.B(net1144),
    .A(net528),
    .X(_2050_));
 sg13g2_or2_1 _5288_ (.X(_2051_),
    .B(_2050_),
    .A(_2048_));
 sg13g2_nand2_1 _5289_ (.Y(_2052_),
    .A(net496),
    .B(_2051_));
 sg13g2_a21oi_1 _5290_ (.A1(_2048_),
    .A2(_2050_),
    .Y(_0294_),
    .B1(_2052_));
 sg13g2_xor2_1 _5291_ (.B(net1259),
    .A(net528),
    .X(_2053_));
 sg13g2_a21oi_1 _5292_ (.A1(_2049_),
    .A2(_2051_),
    .Y(_2054_),
    .B1(_2053_));
 sg13g2_and3_1 _5293_ (.X(_2055_),
    .A(_2049_),
    .B(_2051_),
    .C(_2053_));
 sg13g2_nor3_1 _5294_ (.A(net435),
    .B(_2054_),
    .C(_2055_),
    .Y(_0295_));
 sg13g2_nor2_1 _5295_ (.A(_2051_),
    .B(_2053_),
    .Y(_2056_));
 sg13g2_o21ai_1 _5296_ (.B1(_2049_),
    .Y(_2057_),
    .A1(net528),
    .A2(_0572_));
 sg13g2_nor2_1 _5297_ (.A(_2056_),
    .B(_2057_),
    .Y(_2058_));
 sg13g2_nand2_1 _5298_ (.Y(_2059_),
    .A(net415),
    .B(net1313));
 sg13g2_xor2_1 _5299_ (.B(net1313),
    .A(net529),
    .X(_2060_));
 sg13g2_or2_1 _5300_ (.X(_2061_),
    .B(_2060_),
    .A(_2058_));
 sg13g2_nand2_1 _5301_ (.Y(_2062_),
    .A(net497),
    .B(_2061_));
 sg13g2_a21oi_1 _5302_ (.A1(_2058_),
    .A2(_2060_),
    .Y(_0296_),
    .B1(_2062_));
 sg13g2_xor2_1 _5303_ (.B(net1268),
    .A(net529),
    .X(_2063_));
 sg13g2_and3_1 _5304_ (.X(_2064_),
    .A(_2059_),
    .B(_2061_),
    .C(_2063_));
 sg13g2_a21oi_1 _5305_ (.A1(_2059_),
    .A2(_2061_),
    .Y(_2065_),
    .B1(_2063_));
 sg13g2_nor3_1 _5306_ (.A(net435),
    .B(_2064_),
    .C(net1269),
    .Y(_0297_));
 sg13g2_nor2_1 _5307_ (.A(_2060_),
    .B(_2063_),
    .Y(_2066_));
 sg13g2_nand2b_1 _5308_ (.Y(_2067_),
    .B(_2059_),
    .A_N(_2057_));
 sg13g2_a221oi_1 _5309_ (.B2(_2066_),
    .C1(_2067_),
    .B1(_2056_),
    .A1(net415),
    .Y(_2068_),
    .A2(net1268));
 sg13g2_xor2_1 _5310_ (.B(net837),
    .A(net529),
    .X(_2069_));
 sg13g2_o21ai_1 _5311_ (.B1(net496),
    .Y(_2070_),
    .A1(_2068_),
    .A2(_2069_));
 sg13g2_a21oi_1 _5312_ (.A1(_2068_),
    .A2(_2069_),
    .Y(_0298_),
    .B1(_2070_));
 sg13g2_a21oi_1 _5313_ (.A1(_0564_),
    .A2(net837),
    .Y(_0299_),
    .B1(_2070_));
 sg13g2_nand2_1 _5314_ (.Y(_2071_),
    .A(net970),
    .B(net1008));
 sg13g2_o21ai_1 _5315_ (.B1(net477),
    .Y(_2072_),
    .A1(net970),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[0] ));
 sg13g2_nor2b_1 _5316_ (.A(net971),
    .B_N(_2071_),
    .Y(_0300_));
 sg13g2_nor2b_1 _5317_ (.A(net521),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[0] ),
    .Y(_2073_));
 sg13g2_xnor2_1 _5318_ (.Y(_2074_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[1] ),
    .B(_2073_));
 sg13g2_or2_1 _5319_ (.X(_2075_),
    .B(_2074_),
    .A(_0554_));
 sg13g2_xnor2_1 _5320_ (.Y(_2076_),
    .A(_0554_),
    .B(_2074_));
 sg13g2_o21ai_1 _5321_ (.B1(net477),
    .Y(_2077_),
    .A1(_2071_),
    .A2(_2076_));
 sg13g2_a21oi_1 _5322_ (.A1(_2071_),
    .A2(_2076_),
    .Y(_0301_),
    .B1(_2077_));
 sg13g2_o21ai_1 _5323_ (.B1(_2075_),
    .Y(_2078_),
    .A1(_2071_),
    .A2(_2076_));
 sg13g2_o21ai_1 _5324_ (.B1(net418),
    .Y(_2079_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[0] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[1] ));
 sg13g2_xnor2_1 _5325_ (.Y(_2080_),
    .A(_0555_),
    .B(_2079_));
 sg13g2_nor2_1 _5326_ (.A(_0556_),
    .B(_2080_),
    .Y(_2081_));
 sg13g2_nand2_1 _5327_ (.Y(_2082_),
    .A(_0556_),
    .B(_2080_));
 sg13g2_nand2b_1 _5328_ (.Y(_2083_),
    .B(_2082_),
    .A_N(_2081_));
 sg13g2_nor2b_1 _5329_ (.A(_2078_),
    .B_N(_2083_),
    .Y(_2084_));
 sg13g2_nor2b_1 _5330_ (.A(_2083_),
    .B_N(_2078_),
    .Y(_2085_));
 sg13g2_nor3_1 _5331_ (.A(net429),
    .B(_2084_),
    .C(_2085_),
    .Y(_0302_));
 sg13g2_a21oi_1 _5332_ (.A1(_2078_),
    .A2(_2082_),
    .Y(_2086_),
    .B1(_2081_));
 sg13g2_o21ai_1 _5333_ (.B1(_2079_),
    .Y(_2087_),
    .A1(net521),
    .A2(_0555_));
 sg13g2_xor2_1 _5334_ (.B(_2087_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[3] ),
    .X(_2088_));
 sg13g2_nand2_1 _5335_ (.Y(_2089_),
    .A(net1255),
    .B(_2088_));
 sg13g2_xnor2_1 _5336_ (.Y(_2090_),
    .A(net1255),
    .B(_2088_));
 sg13g2_o21ai_1 _5337_ (.B1(net477),
    .Y(_2091_),
    .A1(_2086_),
    .A2(_2090_));
 sg13g2_a21oi_1 _5338_ (.A1(_2086_),
    .A2(net1256),
    .Y(_0303_),
    .B1(_2091_));
 sg13g2_o21ai_1 _5339_ (.B1(_2089_),
    .Y(_2092_),
    .A1(_2086_),
    .A2(_2090_));
 sg13g2_nor2b_1 _5340_ (.A(net521),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[3] ),
    .Y(_2093_));
 sg13g2_nor3_2 _5341_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[4] ),
    .B(_2087_),
    .C(_2093_),
    .Y(_2094_));
 sg13g2_inv_1 _5342_ (.Y(_2095_),
    .A(_2094_));
 sg13g2_o21ai_1 _5343_ (.B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[4] ),
    .Y(_2096_),
    .A1(_2087_),
    .A2(_2093_));
 sg13g2_nor2b_1 _5344_ (.A(_2094_),
    .B_N(_2096_),
    .Y(_2097_));
 sg13g2_and2_1 _5345_ (.A(net1505),
    .B(_2097_),
    .X(_2098_));
 sg13g2_or2_1 _5346_ (.X(_2099_),
    .B(_2097_),
    .A(net1505));
 sg13g2_nor2b_1 _5347_ (.A(_2098_),
    .B_N(_2099_),
    .Y(_2100_));
 sg13g2_nor2_1 _5348_ (.A(_2092_),
    .B(_2100_),
    .Y(_2101_));
 sg13g2_a21oi_1 _5349_ (.A1(_2092_),
    .A2(_2100_),
    .Y(_2102_),
    .B1(net429));
 sg13g2_nor2b_1 _5350_ (.A(_2101_),
    .B_N(_2102_),
    .Y(_0304_));
 sg13g2_a21oi_1 _5351_ (.A1(_2092_),
    .A2(_2099_),
    .Y(_2103_),
    .B1(_2098_));
 sg13g2_nor2_1 _5352_ (.A(net521),
    .B(_2094_),
    .Y(_2104_));
 sg13g2_xnor2_1 _5353_ (.Y(_2105_),
    .A(_0557_),
    .B(_2104_));
 sg13g2_nand2_1 _5354_ (.Y(_2106_),
    .A(net1417),
    .B(_2105_));
 sg13g2_xnor2_1 _5355_ (.Y(_2107_),
    .A(net1417),
    .B(_2105_));
 sg13g2_o21ai_1 _5356_ (.B1(net478),
    .Y(_2108_),
    .A1(_2103_),
    .A2(_2107_));
 sg13g2_a21oi_1 _5357_ (.A1(_2103_),
    .A2(_2107_),
    .Y(_0305_),
    .B1(_2108_));
 sg13g2_o21ai_1 _5358_ (.B1(_2106_),
    .Y(_2109_),
    .A1(_2103_),
    .A2(_2107_));
 sg13g2_a21oi_1 _5359_ (.A1(_0557_),
    .A2(_2094_),
    .Y(_2110_),
    .B1(net522));
 sg13g2_xor2_1 _5360_ (.B(_2110_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[6] ),
    .X(_2111_));
 sg13g2_and2_1 _5361_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][6] ),
    .B(_2111_),
    .X(_2112_));
 sg13g2_xnor2_1 _5362_ (.Y(_2113_),
    .A(net1541),
    .B(_2111_));
 sg13g2_inv_1 _5363_ (.Y(_2114_),
    .A(_2113_));
 sg13g2_nor2_1 _5364_ (.A(_2109_),
    .B(_2114_),
    .Y(_2115_));
 sg13g2_and2_1 _5365_ (.A(_2109_),
    .B(_2114_),
    .X(_2116_));
 sg13g2_nor3_1 _5366_ (.A(net429),
    .B(_2115_),
    .C(_2116_),
    .Y(_0306_));
 sg13g2_a21oi_1 _5367_ (.A1(_2109_),
    .A2(_2114_),
    .Y(_2117_),
    .B1(_2112_));
 sg13g2_nor3_1 _5368_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[5] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[6] ),
    .C(_2095_),
    .Y(_2118_));
 sg13g2_nor2_1 _5369_ (.A(net522),
    .B(_2118_),
    .Y(_2119_));
 sg13g2_xnor2_1 _5370_ (.Y(_2120_),
    .A(_0559_),
    .B(_2119_));
 sg13g2_nand2_1 _5371_ (.Y(_2121_),
    .A(net1444),
    .B(_2120_));
 sg13g2_xnor2_1 _5372_ (.Y(_2122_),
    .A(net1444),
    .B(_2120_));
 sg13g2_o21ai_1 _5373_ (.B1(net477),
    .Y(_2123_),
    .A1(_2117_),
    .A2(_2122_));
 sg13g2_a21oi_1 _5374_ (.A1(_2117_),
    .A2(_2122_),
    .Y(_0307_),
    .B1(_2123_));
 sg13g2_o21ai_1 _5375_ (.B1(_2121_),
    .Y(_2124_),
    .A1(_2117_),
    .A2(_2122_));
 sg13g2_a21oi_1 _5376_ (.A1(_0559_),
    .A2(_2118_),
    .Y(_2125_),
    .B1(net522));
 sg13g2_xor2_1 _5377_ (.B(_2125_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[10] ),
    .X(_2126_));
 sg13g2_and2_1 _5378_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][8] ),
    .B(_2126_),
    .X(_2127_));
 sg13g2_xnor2_1 _5379_ (.Y(_2128_),
    .A(_0560_),
    .B(_2126_));
 sg13g2_or2_1 _5380_ (.X(_2129_),
    .B(_2128_),
    .A(_2124_));
 sg13g2_nand2_1 _5381_ (.Y(_2130_),
    .A(_2124_),
    .B(_2128_));
 sg13g2_and3_1 _5382_ (.X(_0308_),
    .A(net478),
    .B(_2129_),
    .C(_2130_));
 sg13g2_nand2b_1 _5383_ (.Y(_2131_),
    .B(_2130_),
    .A_N(_2127_));
 sg13g2_mux2_1 _5384_ (.A0(_2125_),
    .A1(net522),
    .S(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[10] ),
    .X(_2132_));
 sg13g2_nor2_1 _5385_ (.A(net1390),
    .B(_2132_),
    .Y(_2133_));
 sg13g2_xor2_1 _5386_ (.B(_2132_),
    .A(net1390),
    .X(_2134_));
 sg13g2_o21ai_1 _5387_ (.B1(net478),
    .Y(_2135_),
    .A1(_2131_),
    .A2(_2134_));
 sg13g2_a21oi_1 _5388_ (.A1(_2131_),
    .A2(_2134_),
    .Y(_0309_),
    .B1(_2135_));
 sg13g2_and2_1 _5389_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][10] ),
    .B(_2132_),
    .X(_2136_));
 sg13g2_xor2_1 _5390_ (.B(_2132_),
    .A(net1479),
    .X(_2137_));
 sg13g2_a221oi_1 _5391_ (.B2(net1390),
    .C1(_2127_),
    .B1(_2132_),
    .A1(_2124_),
    .Y(_2138_),
    .A2(_2128_));
 sg13g2_nor2_1 _5392_ (.A(_2133_),
    .B(_2138_),
    .Y(_2139_));
 sg13g2_o21ai_1 _5393_ (.B1(net477),
    .Y(_2140_),
    .A1(_2137_),
    .A2(_2139_));
 sg13g2_a21oi_1 _5394_ (.A1(_2137_),
    .A2(_2139_),
    .Y(_0310_),
    .B1(_2140_));
 sg13g2_a21oi_1 _5395_ (.A1(_2137_),
    .A2(_2139_),
    .Y(_2141_),
    .B1(_2136_));
 sg13g2_nor2_1 _5396_ (.A(net1386),
    .B(_2132_),
    .Y(_2142_));
 sg13g2_nand2_1 _5397_ (.Y(_2143_),
    .A(net1386),
    .B(_2132_));
 sg13g2_nand2b_1 _5398_ (.Y(_2144_),
    .B(_2143_),
    .A_N(_2142_));
 sg13g2_o21ai_1 _5399_ (.B1(net478),
    .Y(_2145_),
    .A1(_2141_),
    .A2(_2144_));
 sg13g2_a21oi_1 _5400_ (.A1(_2141_),
    .A2(_2144_),
    .Y(_0311_),
    .B1(_2145_));
 sg13g2_o21ai_1 _5401_ (.B1(_2143_),
    .Y(_2146_),
    .A1(_2141_),
    .A2(_2142_));
 sg13g2_xor2_1 _5402_ (.B(_2132_),
    .A(net1233),
    .X(_2147_));
 sg13g2_o21ai_1 _5403_ (.B1(net479),
    .Y(_2148_),
    .A1(_2146_),
    .A2(_2147_));
 sg13g2_a21oi_1 _5404_ (.A1(_2146_),
    .A2(_2147_),
    .Y(_0312_),
    .B1(_2148_));
 sg13g2_nor2b_1 _5405_ (.A(net1054),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][4] ),
    .Y(_2149_));
 sg13g2_xnor2_1 _5406_ (.Y(_2150_),
    .A(net1054),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][4] ));
 sg13g2_nor2_1 _5407_ (.A(net439),
    .B(net1055),
    .Y(_0313_));
 sg13g2_nor2b_1 _5408_ (.A(net521),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][4] ),
    .Y(_2151_));
 sg13g2_xnor2_1 _5409_ (.Y(_2152_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][5] ),
    .B(_2151_));
 sg13g2_nand2_1 _5410_ (.Y(_2153_),
    .A(net1304),
    .B(_2152_));
 sg13g2_xnor2_1 _5411_ (.Y(_2154_),
    .A(net1304),
    .B(_2152_));
 sg13g2_o21ai_1 _5412_ (.B1(net477),
    .Y(_2155_),
    .A1(_2149_),
    .A2(_2154_));
 sg13g2_a21oi_1 _5413_ (.A1(_2149_),
    .A2(_2154_),
    .Y(_0314_),
    .B1(_2155_));
 sg13g2_o21ai_1 _5414_ (.B1(_2153_),
    .Y(_2156_),
    .A1(_2149_),
    .A2(_2154_));
 sg13g2_nor2_1 _5415_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][4] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][5] ),
    .Y(_2157_));
 sg13g2_nor2_1 _5416_ (.A(net521),
    .B(_2157_),
    .Y(_2158_));
 sg13g2_xnor2_1 _5417_ (.Y(_2159_),
    .A(_0558_),
    .B(_2158_));
 sg13g2_nor2b_1 _5418_ (.A(_2159_),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[4][2] ),
    .Y(_2160_));
 sg13g2_xnor2_1 _5419_ (.Y(_2161_),
    .A(net1379),
    .B(_2159_));
 sg13g2_nor2_1 _5420_ (.A(_2156_),
    .B(_2161_),
    .Y(_2162_));
 sg13g2_a21oi_1 _5421_ (.A1(_2156_),
    .A2(_2161_),
    .Y(_2163_),
    .B1(net429));
 sg13g2_nor2b_1 _5422_ (.A(_2162_),
    .B_N(_2163_),
    .Y(_0315_));
 sg13g2_a21oi_1 _5423_ (.A1(_2156_),
    .A2(_2161_),
    .Y(_2164_),
    .B1(_2160_));
 sg13g2_a21oi_1 _5424_ (.A1(_0558_),
    .A2(_2157_),
    .Y(_2165_),
    .B1(net521));
 sg13g2_xnor2_1 _5425_ (.Y(_2166_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][7] ),
    .B(_2165_));
 sg13g2_nand2_1 _5426_ (.Y(_2167_),
    .A(net1367),
    .B(_2166_));
 sg13g2_xor2_1 _5427_ (.B(_2166_),
    .A(net1367),
    .X(_2168_));
 sg13g2_inv_1 _5428_ (.Y(_2169_),
    .A(_2168_));
 sg13g2_o21ai_1 _5429_ (.B1(net477),
    .Y(_2170_),
    .A1(_2164_),
    .A2(_2169_));
 sg13g2_a21oi_1 _5430_ (.A1(_2164_),
    .A2(_2169_),
    .Y(_0316_),
    .B1(_2170_));
 sg13g2_o21ai_1 _5431_ (.B1(_2167_),
    .Y(_2171_),
    .A1(_2164_),
    .A2(_2169_));
 sg13g2_a21oi_1 _5432_ (.A1(net418),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][7] ),
    .Y(_2172_),
    .B1(_2165_));
 sg13g2_xnor2_1 _5433_ (.Y(_2173_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][8] ),
    .B(_2172_));
 sg13g2_nor2b_1 _5434_ (.A(_2173_),
    .B_N(net1008),
    .Y(_2174_));
 sg13g2_xnor2_1 _5435_ (.Y(_2175_),
    .A(net1008),
    .B(_2173_));
 sg13g2_nor2_1 _5436_ (.A(_2171_),
    .B(_2175_),
    .Y(_2176_));
 sg13g2_a21oi_1 _5437_ (.A1(_2171_),
    .A2(_2175_),
    .Y(_2177_),
    .B1(net429));
 sg13g2_nor2b_1 _5438_ (.A(_2176_),
    .B_N(_2177_),
    .Y(_0317_));
 sg13g2_a21oi_1 _5439_ (.A1(_2171_),
    .A2(_2175_),
    .Y(_2178_),
    .B1(_2174_));
 sg13g2_a21oi_1 _5440_ (.A1(_0560_),
    .A2(_2172_),
    .Y(_2179_),
    .B1(net521));
 sg13g2_xnor2_1 _5441_ (.Y(_2180_),
    .A(net1570),
    .B(_2179_));
 sg13g2_nand2_1 _5442_ (.Y(_2181_),
    .A(net1317),
    .B(_2180_));
 sg13g2_nor2_1 _5443_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[1] ),
    .B(_2180_),
    .Y(_2182_));
 sg13g2_xor2_1 _5444_ (.B(_2180_),
    .A(net1317),
    .X(_2183_));
 sg13g2_nor2b_1 _5445_ (.A(_2183_),
    .B_N(_2178_),
    .Y(_2184_));
 sg13g2_nor2b_1 _5446_ (.A(_2178_),
    .B_N(_2183_),
    .Y(_2185_));
 sg13g2_nor3_1 _5447_ (.A(net429),
    .B(_2184_),
    .C(_2185_),
    .Y(_0318_));
 sg13g2_o21ai_1 _5448_ (.B1(_2181_),
    .Y(_2186_),
    .A1(_2178_),
    .A2(_2182_));
 sg13g2_a21o_1 _5449_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][9] ),
    .A1(net418),
    .B1(_2179_),
    .X(_2187_));
 sg13g2_xnor2_1 _5450_ (.Y(_2188_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][10] ),
    .B(_2187_));
 sg13g2_and2_1 _5451_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[2] ),
    .B(_2188_),
    .X(_2189_));
 sg13g2_xnor2_1 _5452_ (.Y(_2190_),
    .A(_0555_),
    .B(_2188_));
 sg13g2_or2_1 _5453_ (.X(_2191_),
    .B(_2190_),
    .A(_2186_));
 sg13g2_a21oi_1 _5454_ (.A1(_2186_),
    .A2(_2190_),
    .Y(_2192_),
    .B1(net429));
 sg13g2_and2_1 _5455_ (.A(_2191_),
    .B(_2192_),
    .X(_0319_));
 sg13g2_a21oi_1 _5456_ (.A1(_2186_),
    .A2(_2190_),
    .Y(_2193_),
    .B1(_2189_));
 sg13g2_a21o_1 _5457_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][10] ),
    .A1(net418),
    .B1(_2187_),
    .X(_2194_));
 sg13g2_xnor2_1 _5458_ (.Y(_2195_),
    .A(net1386),
    .B(_2194_));
 sg13g2_nand2_1 _5459_ (.Y(_2196_),
    .A(net1388),
    .B(_2195_));
 sg13g2_xnor2_1 _5460_ (.Y(_2197_),
    .A(net1388),
    .B(_2195_));
 sg13g2_o21ai_1 _5461_ (.B1(net477),
    .Y(_2198_),
    .A1(_2193_),
    .A2(_2197_));
 sg13g2_a21oi_1 _5462_ (.A1(_2193_),
    .A2(_2197_),
    .Y(_0320_),
    .B1(_2198_));
 sg13g2_o21ai_1 _5463_ (.B1(_2196_),
    .Y(_2199_),
    .A1(_2193_),
    .A2(_2197_));
 sg13g2_a21o_1 _5464_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][11] ),
    .A1(net418),
    .B1(_2194_),
    .X(_2200_));
 sg13g2_xnor2_1 _5465_ (.Y(_2201_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][12] ),
    .B(_2200_));
 sg13g2_nand2_1 _5466_ (.Y(_2202_),
    .A(net1502),
    .B(_2201_));
 sg13g2_xnor2_1 _5467_ (.Y(_2203_),
    .A(net1502),
    .B(_2201_));
 sg13g2_nand2b_1 _5468_ (.Y(_2204_),
    .B(_2203_),
    .A_N(_2199_));
 sg13g2_nand2b_1 _5469_ (.Y(_2205_),
    .B(_2199_),
    .A_N(_2203_));
 sg13g2_and3_1 _5470_ (.X(_0321_),
    .A(net479),
    .B(_2204_),
    .C(_2205_));
 sg13g2_mux2_1 _5471_ (.A0(_2200_),
    .A1(net522),
    .S(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][12] ),
    .X(_2206_));
 sg13g2_inv_1 _5472_ (.Y(_2207_),
    .A(_2206_));
 sg13g2_xnor2_1 _5473_ (.Y(_2208_),
    .A(_0557_),
    .B(_2206_));
 sg13g2_a21oi_1 _5474_ (.A1(_2202_),
    .A2(_2205_),
    .Y(_2209_),
    .B1(_2208_));
 sg13g2_and3_1 _5475_ (.X(_2210_),
    .A(_2202_),
    .B(_2205_),
    .C(_2208_));
 sg13g2_nor3_1 _5476_ (.A(net430),
    .B(_2209_),
    .C(_2210_),
    .Y(_0322_));
 sg13g2_nand2_1 _5477_ (.Y(_2211_),
    .A(net1483),
    .B(_2207_));
 sg13g2_xor2_1 _5478_ (.B(_2206_),
    .A(net1483),
    .X(_2212_));
 sg13g2_or2_1 _5479_ (.X(_2213_),
    .B(_2208_),
    .A(_2205_));
 sg13g2_o21ai_1 _5480_ (.B1(_2202_),
    .Y(_2214_),
    .A1(_0557_),
    .A2(_2206_));
 sg13g2_inv_1 _5481_ (.Y(_2215_),
    .A(_2214_));
 sg13g2_nand3_1 _5482_ (.B(_2213_),
    .C(_2215_),
    .A(_2212_),
    .Y(_2216_));
 sg13g2_a21o_1 _5483_ (.A2(_2215_),
    .A1(_2213_),
    .B1(_2212_),
    .X(_2217_));
 sg13g2_and3_1 _5484_ (.X(_0323_),
    .A(net479),
    .B(_2216_),
    .C(_2217_));
 sg13g2_xnor2_1 _5485_ (.Y(_2218_),
    .A(_0559_),
    .B(_2206_));
 sg13g2_and3_1 _5486_ (.X(_2219_),
    .A(_2211_),
    .B(_2217_),
    .C(_2218_));
 sg13g2_a21oi_1 _5487_ (.A1(_2211_),
    .A2(_2217_),
    .Y(_2220_),
    .B1(_2218_));
 sg13g2_nor3_1 _5488_ (.A(net430),
    .B(_2219_),
    .C(net1484),
    .Y(_0324_));
 sg13g2_nor3_1 _5489_ (.A(_2212_),
    .B(_2213_),
    .C(_2218_),
    .Y(_2221_));
 sg13g2_o21ai_1 _5490_ (.B1(_2211_),
    .Y(_2222_),
    .A1(_0559_),
    .A2(_2206_));
 sg13g2_nor3_1 _5491_ (.A(_2214_),
    .B(_2221_),
    .C(_2222_),
    .Y(_2223_));
 sg13g2_xor2_1 _5492_ (.B(_2206_),
    .A(net1285),
    .X(_2224_));
 sg13g2_o21ai_1 _5493_ (.B1(net479),
    .Y(_2225_),
    .A1(_2223_),
    .A2(_2224_));
 sg13g2_a21oi_1 _5494_ (.A1(_2223_),
    .A2(_2224_),
    .Y(_0325_),
    .B1(_2225_));
 sg13g2_nor2_1 _5495_ (.A(net852),
    .B(net432),
    .Y(_0326_));
 sg13g2_nor2b_1 _5496_ (.A(net524),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][1] ),
    .Y(_2226_));
 sg13g2_xnor2_1 _5497_ (.Y(_2227_),
    .A(net524),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][1] ));
 sg13g2_o21ai_1 _5498_ (.B1(net482),
    .Y(_2228_),
    .A1(net852),
    .A2(_2227_));
 sg13g2_a21oi_1 _5499_ (.A1(net852),
    .A2(_2227_),
    .Y(_0327_),
    .B1(_2228_));
 sg13g2_a21oi_1 _5500_ (.A1(net852),
    .A2(_2227_),
    .Y(_2229_),
    .B1(_2226_));
 sg13g2_nand2_1 _5501_ (.Y(_2230_),
    .A(net418),
    .B(net1074));
 sg13g2_xor2_1 _5502_ (.B(net1074),
    .A(net524),
    .X(_2231_));
 sg13g2_or2_1 _5503_ (.X(_2232_),
    .B(_2231_),
    .A(_2229_));
 sg13g2_nand2_1 _5504_ (.Y(_2233_),
    .A(net481),
    .B(_2232_));
 sg13g2_a21oi_1 _5505_ (.A1(_2229_),
    .A2(_2231_),
    .Y(_0328_),
    .B1(_2233_));
 sg13g2_xnor2_1 _5506_ (.Y(_2234_),
    .A(net524),
    .B(net1089));
 sg13g2_nand3_1 _5507_ (.B(_2232_),
    .C(_2234_),
    .A(_2230_),
    .Y(_2235_));
 sg13g2_a21o_1 _5508_ (.A2(_2232_),
    .A1(_2230_),
    .B1(_2234_),
    .X(_2236_));
 sg13g2_inv_1 _5509_ (.Y(_2237_),
    .A(_2236_));
 sg13g2_and3_1 _5510_ (.X(_0329_),
    .A(net481),
    .B(_2235_),
    .C(_2236_));
 sg13g2_a21oi_1 _5511_ (.A1(net524),
    .A2(net1089),
    .Y(_2238_),
    .B1(_2237_));
 sg13g2_nand2_1 _5512_ (.Y(_2239_),
    .A(net418),
    .B(net1358));
 sg13g2_xor2_1 _5513_ (.B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][4] ),
    .A(net523),
    .X(_2240_));
 sg13g2_or2_1 _5514_ (.X(_2241_),
    .B(_2240_),
    .A(_2238_));
 sg13g2_nand2_1 _5515_ (.Y(_2242_),
    .A(net481),
    .B(_2241_));
 sg13g2_a21oi_1 _5516_ (.A1(_2238_),
    .A2(_2240_),
    .Y(_0330_),
    .B1(_2242_));
 sg13g2_and2_1 _5517_ (.A(_2239_),
    .B(_2241_),
    .X(_2243_));
 sg13g2_nor2_1 _5518_ (.A(net523),
    .B(net1563),
    .Y(_2244_));
 sg13g2_and2_1 _5519_ (.A(net523),
    .B(net1563),
    .X(_2245_));
 sg13g2_or2_1 _5520_ (.X(_2246_),
    .B(_2245_),
    .A(_2244_));
 sg13g2_o21ai_1 _5521_ (.B1(net481),
    .Y(_2247_),
    .A1(_2243_),
    .A2(_2246_));
 sg13g2_a21oi_1 _5522_ (.A1(_2243_),
    .A2(_2246_),
    .Y(_0331_),
    .B1(_2247_));
 sg13g2_xnor2_1 _5523_ (.Y(_2248_),
    .A(net523),
    .B(net1506));
 sg13g2_nor2_1 _5524_ (.A(_2243_),
    .B(_2244_),
    .Y(_2249_));
 sg13g2_or3_1 _5525_ (.A(_2245_),
    .B(_2248_),
    .C(_2249_),
    .X(_2250_));
 sg13g2_o21ai_1 _5526_ (.B1(_2248_),
    .Y(_2251_),
    .A1(_2245_),
    .A2(_2249_));
 sg13g2_and3_1 _5527_ (.X(_0332_),
    .A(net481),
    .B(_2250_),
    .C(_2251_));
 sg13g2_o21ai_1 _5528_ (.B1(_2251_),
    .Y(_2252_),
    .A1(net523),
    .A2(_0561_));
 sg13g2_xnor2_1 _5529_ (.Y(_2253_),
    .A(net523),
    .B(net1156));
 sg13g2_o21ai_1 _5530_ (.B1(net481),
    .Y(_2254_),
    .A1(_2252_),
    .A2(_2253_));
 sg13g2_a21oi_1 _5531_ (.A1(_2252_),
    .A2(_2253_),
    .Y(_0333_),
    .B1(_2254_));
 sg13g2_nand2b_1 _5532_ (.Y(_2255_),
    .B(_2253_),
    .A_N(_2251_));
 sg13g2_o21ai_1 _5533_ (.B1(net418),
    .Y(_2256_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][6] ),
    .A2(net1156));
 sg13g2_and2_1 _5534_ (.A(_2255_),
    .B(net1507),
    .X(_2257_));
 sg13g2_xor2_1 _5535_ (.B(net1124),
    .A(net523),
    .X(_2258_));
 sg13g2_and2_1 _5536_ (.A(_2257_),
    .B(_2258_),
    .X(_2259_));
 sg13g2_nor2_1 _5537_ (.A(_2257_),
    .B(_2258_),
    .Y(_2260_));
 sg13g2_nor3_1 _5538_ (.A(net432),
    .B(_2259_),
    .C(_2260_),
    .Y(_0334_));
 sg13g2_a21o_1 _5539_ (.A2(net1124),
    .A1(_0553_),
    .B1(_2260_),
    .X(_2261_));
 sg13g2_nor2b_1 _5540_ (.A(net525),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][9] ),
    .Y(_2262_));
 sg13g2_xnor2_1 _5541_ (.Y(_2263_),
    .A(net525),
    .B(net1171));
 sg13g2_o21ai_1 _5542_ (.B1(net476),
    .Y(_2264_),
    .A1(_2261_),
    .A2(_2263_));
 sg13g2_a21oi_1 _5543_ (.A1(_2261_),
    .A2(net1172),
    .Y(_0335_),
    .B1(_2264_));
 sg13g2_a221oi_1 _5544_ (.B2(_2263_),
    .C1(_2262_),
    .B1(_2260_),
    .A1(_0553_),
    .Y(_2265_),
    .A2(net1124));
 sg13g2_xor2_1 _5545_ (.B(net811),
    .A(net525),
    .X(_2266_));
 sg13g2_o21ai_1 _5546_ (.B1(net479),
    .Y(_2267_),
    .A1(net1125),
    .A2(_2266_));
 sg13g2_a21oi_1 _5547_ (.A1(net1125),
    .A2(_2266_),
    .Y(_0336_),
    .B1(_2267_));
 sg13g2_a21oi_1 _5548_ (.A1(_0553_),
    .A2(net811),
    .Y(_0337_),
    .B1(_2267_));
 sg13g2_and2_1 _5549_ (.A(net933),
    .B(net1230),
    .X(_2268_));
 sg13g2_o21ai_1 _5550_ (.B1(net474),
    .Y(_2269_),
    .A1(net933),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[0] ));
 sg13g2_nor2_1 _5551_ (.A(_2268_),
    .B(net934),
    .Y(_0338_));
 sg13g2_nor2b_1 _5552_ (.A(net515),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[0] ),
    .Y(_2270_));
 sg13g2_xnor2_1 _5553_ (.Y(_2271_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[1] ),
    .B(_2270_));
 sg13g2_nor2_1 _5554_ (.A(_0593_),
    .B(_2271_),
    .Y(_2272_));
 sg13g2_nand2_1 _5555_ (.Y(_2273_),
    .A(_0593_),
    .B(_2271_));
 sg13g2_nor2b_1 _5556_ (.A(_2272_),
    .B_N(_2273_),
    .Y(_2274_));
 sg13g2_nor2_1 _5557_ (.A(_2268_),
    .B(_2274_),
    .Y(_2275_));
 sg13g2_a21oi_1 _5558_ (.A1(_2268_),
    .A2(_2274_),
    .Y(_2276_),
    .B1(net425));
 sg13g2_nor2b_1 _5559_ (.A(net1231),
    .B_N(_2276_),
    .Y(_0339_));
 sg13g2_a21oi_1 _5560_ (.A1(_2268_),
    .A2(_2273_),
    .Y(_2277_),
    .B1(_2272_));
 sg13g2_nor2_1 _5561_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[0] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[1] ),
    .Y(_2278_));
 sg13g2_nor2_1 _5562_ (.A(net515),
    .B(_2278_),
    .Y(_2279_));
 sg13g2_xnor2_1 _5563_ (.Y(_2280_),
    .A(_0594_),
    .B(_2279_));
 sg13g2_nand2_1 _5564_ (.Y(_2281_),
    .A(net1302),
    .B(_2280_));
 sg13g2_xnor2_1 _5565_ (.Y(_2282_),
    .A(net1302),
    .B(_2280_));
 sg13g2_o21ai_1 _5566_ (.B1(net474),
    .Y(_2283_),
    .A1(_2277_),
    .A2(_2282_));
 sg13g2_a21oi_1 _5567_ (.A1(_2277_),
    .A2(_2282_),
    .Y(_0340_),
    .B1(_2283_));
 sg13g2_o21ai_1 _5568_ (.B1(_2281_),
    .Y(_2284_),
    .A1(_2277_),
    .A2(_2282_));
 sg13g2_a21oi_1 _5569_ (.A1(_0594_),
    .A2(_2278_),
    .Y(_2285_),
    .B1(net515));
 sg13g2_nor2_1 _5570_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[3] ),
    .B(_2285_),
    .Y(_2286_));
 sg13g2_xor2_1 _5571_ (.B(_2285_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[3] ),
    .X(_2287_));
 sg13g2_nand2_1 _5572_ (.Y(_2288_),
    .A(net1384),
    .B(_2287_));
 sg13g2_inv_1 _5573_ (.Y(_2289_),
    .A(_2288_));
 sg13g2_xnor2_1 _5574_ (.Y(_2290_),
    .A(net1384),
    .B(_2287_));
 sg13g2_inv_1 _5575_ (.Y(_2291_),
    .A(net1385));
 sg13g2_o21ai_1 _5576_ (.B1(net474),
    .Y(_2292_),
    .A1(_2284_),
    .A2(_2291_));
 sg13g2_a21oi_1 _5577_ (.A1(_2284_),
    .A2(_2291_),
    .Y(_0341_),
    .B1(_2292_));
 sg13g2_a21oi_1 _5578_ (.A1(_2284_),
    .A2(_2291_),
    .Y(_2293_),
    .B1(_2289_));
 sg13g2_nor3_1 _5579_ (.A(net515),
    .B(_0595_),
    .C(_2286_),
    .Y(_2294_));
 sg13g2_o21ai_1 _5580_ (.B1(_0595_),
    .Y(_2295_),
    .A1(net515),
    .A2(_2286_));
 sg13g2_nor2b_1 _5581_ (.A(_2294_),
    .B_N(_2295_),
    .Y(_2296_));
 sg13g2_nand2_1 _5582_ (.Y(_2297_),
    .A(net1415),
    .B(_2296_));
 sg13g2_xnor2_1 _5583_ (.Y(_2298_),
    .A(net1415),
    .B(_2296_));
 sg13g2_o21ai_1 _5584_ (.B1(net474),
    .Y(_2299_),
    .A1(_2293_),
    .A2(_2298_));
 sg13g2_a21oi_1 _5585_ (.A1(_2293_),
    .A2(_2298_),
    .Y(_0342_),
    .B1(_2299_));
 sg13g2_o21ai_1 _5586_ (.B1(_2297_),
    .Y(_2300_),
    .A1(_2293_),
    .A2(_2298_));
 sg13g2_a21oi_1 _5587_ (.A1(_0595_),
    .A2(_2286_),
    .Y(_2301_),
    .B1(net516));
 sg13g2_xor2_1 _5588_ (.B(_2301_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[5] ),
    .X(_2302_));
 sg13g2_and2_1 _5589_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][5] ),
    .B(_2302_),
    .X(_2303_));
 sg13g2_xnor2_1 _5590_ (.Y(_2304_),
    .A(_0596_),
    .B(_2302_));
 sg13g2_o21ai_1 _5591_ (.B1(net474),
    .Y(_2305_),
    .A1(_2300_),
    .A2(_2304_));
 sg13g2_a21oi_1 _5592_ (.A1(_2300_),
    .A2(_2304_),
    .Y(_0343_),
    .B1(_2305_));
 sg13g2_a21oi_1 _5593_ (.A1(_2300_),
    .A2(_2304_),
    .Y(_2306_),
    .B1(_2303_));
 sg13g2_o21ai_1 _5594_ (.B1(net412),
    .Y(_2307_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[5] ),
    .A2(_2295_));
 sg13g2_xnor2_1 _5595_ (.Y(_2308_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[6] ),
    .B(_2307_));
 sg13g2_nand2_1 _5596_ (.Y(_2309_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][6] ),
    .B(_2308_));
 sg13g2_xnor2_1 _5597_ (.Y(_2310_),
    .A(net1412),
    .B(_2308_));
 sg13g2_o21ai_1 _5598_ (.B1(net475),
    .Y(_2311_),
    .A1(_2306_),
    .A2(_2310_));
 sg13g2_a21oi_1 _5599_ (.A1(_2306_),
    .A2(net1413),
    .Y(_0344_),
    .B1(_2311_));
 sg13g2_o21ai_1 _5600_ (.B1(_2309_),
    .Y(_2312_),
    .A1(_2306_),
    .A2(_2310_));
 sg13g2_nor3_1 _5601_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[5] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[6] ),
    .C(_2295_),
    .Y(_2313_));
 sg13g2_nor2_1 _5602_ (.A(net516),
    .B(_2313_),
    .Y(_2314_));
 sg13g2_xor2_1 _5603_ (.B(_2314_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[7] ),
    .X(_2315_));
 sg13g2_and2_1 _5604_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][7] ),
    .B(_2315_),
    .X(_2316_));
 sg13g2_xnor2_1 _5605_ (.Y(_2317_),
    .A(net1401),
    .B(_2315_));
 sg13g2_inv_1 _5606_ (.Y(_2318_),
    .A(net1402));
 sg13g2_o21ai_1 _5607_ (.B1(net475),
    .Y(_2319_),
    .A1(_2312_),
    .A2(_2318_));
 sg13g2_a21oi_1 _5608_ (.A1(_2312_),
    .A2(_2318_),
    .Y(_0345_),
    .B1(_2319_));
 sg13g2_a21o_1 _5609_ (.A2(_2318_),
    .A1(_2312_),
    .B1(_2316_),
    .X(_2320_));
 sg13g2_nor2b_1 _5610_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[7] ),
    .B_N(_2313_),
    .Y(_2321_));
 sg13g2_nor2_1 _5611_ (.A(net516),
    .B(_2321_),
    .Y(_2322_));
 sg13g2_xnor2_1 _5612_ (.Y(_2323_),
    .A(_0597_),
    .B(_2322_));
 sg13g2_and2_1 _5613_ (.A(net1334),
    .B(_2323_),
    .X(_2324_));
 sg13g2_xor2_1 _5614_ (.B(_2323_),
    .A(net1334),
    .X(_2325_));
 sg13g2_nor2_1 _5615_ (.A(_2320_),
    .B(_2325_),
    .Y(_2326_));
 sg13g2_a21oi_1 _5616_ (.A1(_2320_),
    .A2(_2325_),
    .Y(_2327_),
    .B1(net431));
 sg13g2_nor2b_1 _5617_ (.A(net1335),
    .B_N(_2327_),
    .Y(_0346_));
 sg13g2_a21o_1 _5618_ (.A2(_2325_),
    .A1(_2320_),
    .B1(_2324_),
    .X(_2328_));
 sg13g2_a21oi_1 _5619_ (.A1(_0597_),
    .A2(_2321_),
    .Y(_2329_),
    .B1(net516));
 sg13g2_xnor2_1 _5620_ (.Y(_2330_),
    .A(_0598_),
    .B(_2329_));
 sg13g2_and2_1 _5621_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][9] ),
    .B(_2330_),
    .X(_2331_));
 sg13g2_xnor2_1 _5622_ (.Y(_2332_),
    .A(_0599_),
    .B(_2330_));
 sg13g2_o21ai_1 _5623_ (.B1(net474),
    .Y(_2333_),
    .A1(_2328_),
    .A2(_2332_));
 sg13g2_a21oi_1 _5624_ (.A1(_2328_),
    .A2(_2332_),
    .Y(_0347_),
    .B1(_2333_));
 sg13g2_a21o_1 _5625_ (.A2(_2332_),
    .A1(_2328_),
    .B1(_2331_),
    .X(_2334_));
 sg13g2_nor2_1 _5626_ (.A(net412),
    .B(_0598_),
    .Y(_2335_));
 sg13g2_a21oi_2 _5627_ (.B1(_2335_),
    .Y(_2336_),
    .A2(_2329_),
    .A1(_0598_));
 sg13g2_nor2b_1 _5628_ (.A(_2336_),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][10] ),
    .Y(_2337_));
 sg13g2_xnor2_1 _5629_ (.Y(_2338_),
    .A(net1467),
    .B(_2336_));
 sg13g2_nor2_1 _5630_ (.A(_2334_),
    .B(_2338_),
    .Y(_2339_));
 sg13g2_a21oi_1 _5631_ (.A1(_2334_),
    .A2(_2338_),
    .Y(_2340_),
    .B1(net431));
 sg13g2_nor2b_1 _5632_ (.A(net1468),
    .B_N(_2340_),
    .Y(_0348_));
 sg13g2_a21o_1 _5633_ (.A2(_2338_),
    .A1(_2334_),
    .B1(_2337_),
    .X(_2341_));
 sg13g2_nand2b_1 _5634_ (.Y(_2342_),
    .B(_2336_),
    .A_N(net1194));
 sg13g2_nor2b_1 _5635_ (.A(_2336_),
    .B_N(net1194),
    .Y(_2343_));
 sg13g2_xnor2_1 _5636_ (.Y(_2344_),
    .A(net1194),
    .B(_2336_));
 sg13g2_o21ai_1 _5637_ (.B1(net476),
    .Y(_2345_),
    .A1(_2341_),
    .A2(_2344_));
 sg13g2_a21oi_1 _5638_ (.A1(_2341_),
    .A2(_2344_),
    .Y(_0349_),
    .B1(_2345_));
 sg13g2_a21oi_1 _5639_ (.A1(_2341_),
    .A2(_2342_),
    .Y(_2346_),
    .B1(_2343_));
 sg13g2_xor2_1 _5640_ (.B(_2336_),
    .A(net1258),
    .X(_2347_));
 sg13g2_o21ai_1 _5641_ (.B1(net476),
    .Y(_2348_),
    .A1(_2346_),
    .A2(_2347_));
 sg13g2_a21oi_1 _5642_ (.A1(_2346_),
    .A2(_2347_),
    .Y(_0350_),
    .B1(_2348_));
 sg13g2_nor2b_1 _5643_ (.A(net1010),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][3] ),
    .Y(_2349_));
 sg13g2_xnor2_1 _5644_ (.Y(_2350_),
    .A(net1010),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][3] ));
 sg13g2_nor2_1 _5645_ (.A(net431),
    .B(net1011),
    .Y(_0351_));
 sg13g2_nor2b_1 _5646_ (.A(net515),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][3] ),
    .Y(_2351_));
 sg13g2_xnor2_1 _5647_ (.Y(_2352_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][4] ),
    .B(_2351_));
 sg13g2_nand2_1 _5648_ (.Y(_2353_),
    .A(net1240),
    .B(_2352_));
 sg13g2_xnor2_1 _5649_ (.Y(_2354_),
    .A(net1240),
    .B(_2352_));
 sg13g2_o21ai_1 _5650_ (.B1(net474),
    .Y(_2355_),
    .A1(_2349_),
    .A2(_2354_));
 sg13g2_a21oi_1 _5651_ (.A1(_2349_),
    .A2(_2354_),
    .Y(_0352_),
    .B1(_2355_));
 sg13g2_o21ai_1 _5652_ (.B1(_2353_),
    .Y(_2356_),
    .A1(_2349_),
    .A2(_2354_));
 sg13g2_nor2_1 _5653_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][3] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][4] ),
    .Y(_2357_));
 sg13g2_nor2_1 _5654_ (.A(net515),
    .B(_2357_),
    .Y(_2358_));
 sg13g2_xnor2_1 _5655_ (.Y(_2359_),
    .A(_0596_),
    .B(_2358_));
 sg13g2_nor2b_1 _5656_ (.A(_2359_),
    .B_N(net1446),
    .Y(_2360_));
 sg13g2_xnor2_1 _5657_ (.Y(_2361_),
    .A(net1446),
    .B(_2359_));
 sg13g2_nor2_1 _5658_ (.A(_2356_),
    .B(_2361_),
    .Y(_2362_));
 sg13g2_a21oi_1 _5659_ (.A1(_2356_),
    .A2(_2361_),
    .Y(_2363_),
    .B1(net425));
 sg13g2_nor2b_1 _5660_ (.A(_2362_),
    .B_N(_2363_),
    .Y(_0353_));
 sg13g2_a21oi_1 _5661_ (.A1(_2356_),
    .A2(_2361_),
    .Y(_2364_),
    .B1(_2360_));
 sg13g2_a21oi_1 _5662_ (.A1(_0596_),
    .A2(_2357_),
    .Y(_2365_),
    .B1(net515));
 sg13g2_xnor2_1 _5663_ (.Y(_2366_),
    .A(net1412),
    .B(_2365_));
 sg13g2_nand2_1 _5664_ (.Y(_2367_),
    .A(net1230),
    .B(_2366_));
 sg13g2_xor2_1 _5665_ (.B(_2366_),
    .A(net1230),
    .X(_2368_));
 sg13g2_inv_1 _5666_ (.Y(_2369_),
    .A(_2368_));
 sg13g2_o21ai_1 _5667_ (.B1(net474),
    .Y(_2370_),
    .A1(_2364_),
    .A2(_2369_));
 sg13g2_a21oi_1 _5668_ (.A1(_2364_),
    .A2(_2369_),
    .Y(_0354_),
    .B1(_2370_));
 sg13g2_o21ai_1 _5669_ (.B1(_2367_),
    .Y(_2371_),
    .A1(_2364_),
    .A2(_2369_));
 sg13g2_a21oi_1 _5670_ (.A1(net412),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][6] ),
    .Y(_2372_),
    .B1(_2365_));
 sg13g2_nand2b_1 _5671_ (.Y(_2373_),
    .B(_2372_),
    .A_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][7] ));
 sg13g2_xor2_1 _5672_ (.B(_2372_),
    .A(net1401),
    .X(_2374_));
 sg13g2_and2_1 _5673_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[1] ),
    .B(_2374_),
    .X(_2375_));
 sg13g2_xor2_1 _5674_ (.B(_2374_),
    .A(net1443),
    .X(_2376_));
 sg13g2_nor2_1 _5675_ (.A(_2371_),
    .B(_2376_),
    .Y(_2377_));
 sg13g2_a21oi_1 _5676_ (.A1(_2371_),
    .A2(_2376_),
    .Y(_2378_),
    .B1(net431));
 sg13g2_nor2b_1 _5677_ (.A(_2377_),
    .B_N(_2378_),
    .Y(_0355_));
 sg13g2_a21oi_1 _5678_ (.A1(_2371_),
    .A2(_2376_),
    .Y(_2379_),
    .B1(_2375_));
 sg13g2_and2_1 _5679_ (.A(net412),
    .B(_2373_),
    .X(_2380_));
 sg13g2_xnor2_1 _5680_ (.Y(_2381_),
    .A(net1334),
    .B(_2380_));
 sg13g2_nand2_1 _5681_ (.Y(_2382_),
    .A(net1377),
    .B(_2381_));
 sg13g2_xnor2_1 _5682_ (.Y(_2383_),
    .A(net1377),
    .B(_2381_));
 sg13g2_o21ai_1 _5683_ (.B1(net475),
    .Y(_2384_),
    .A1(_2379_),
    .A2(_2383_));
 sg13g2_a21oi_1 _5684_ (.A1(_2379_),
    .A2(_2383_),
    .Y(_0356_),
    .B1(_2384_));
 sg13g2_o21ai_1 _5685_ (.B1(_2382_),
    .Y(_2385_),
    .A1(_2379_),
    .A2(_2383_));
 sg13g2_nor2_1 _5686_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][8] ),
    .B(_2373_),
    .Y(_2386_));
 sg13g2_nor2_1 _5687_ (.A(net516),
    .B(_2386_),
    .Y(_2387_));
 sg13g2_xnor2_1 _5688_ (.Y(_2388_),
    .A(net1482),
    .B(_2387_));
 sg13g2_and2_1 _5689_ (.A(net1456),
    .B(_2388_),
    .X(_2389_));
 sg13g2_xor2_1 _5690_ (.B(_2388_),
    .A(net1456),
    .X(_2390_));
 sg13g2_nor2_1 _5691_ (.A(_2385_),
    .B(_2390_),
    .Y(_2391_));
 sg13g2_a21oi_1 _5692_ (.A1(_2385_),
    .A2(_2390_),
    .Y(_2392_),
    .B1(net431));
 sg13g2_nor2b_1 _5693_ (.A(_2391_),
    .B_N(_2392_),
    .Y(_0357_));
 sg13g2_a21oi_1 _5694_ (.A1(_2385_),
    .A2(_2390_),
    .Y(_2393_),
    .B1(_2389_));
 sg13g2_a21oi_1 _5695_ (.A1(_0599_),
    .A2(_2386_),
    .Y(_2394_),
    .B1(net516));
 sg13g2_xnor2_1 _5696_ (.Y(_2395_),
    .A(net1467),
    .B(_2394_));
 sg13g2_nand2_1 _5697_ (.Y(_2396_),
    .A(net1519),
    .B(_2395_));
 sg13g2_xnor2_1 _5698_ (.Y(_2397_),
    .A(_0595_),
    .B(_2395_));
 sg13g2_inv_1 _5699_ (.Y(_2398_),
    .A(_2397_));
 sg13g2_o21ai_1 _5700_ (.B1(net475),
    .Y(_2399_),
    .A1(_2393_),
    .A2(_2398_));
 sg13g2_a21oi_1 _5701_ (.A1(_2393_),
    .A2(_2398_),
    .Y(_0358_),
    .B1(_2399_));
 sg13g2_o21ai_1 _5702_ (.B1(_2396_),
    .Y(_2400_),
    .A1(_2393_),
    .A2(_2398_));
 sg13g2_a21o_1 _5703_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][10] ),
    .A1(net412),
    .B1(_2394_),
    .X(_2401_));
 sg13g2_xnor2_1 _5704_ (.Y(_2402_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][11] ),
    .B(_2401_));
 sg13g2_and2_1 _5705_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[5] ),
    .B(_2402_),
    .X(_2403_));
 sg13g2_xnor2_1 _5706_ (.Y(_2404_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[5] ),
    .B(_2402_));
 sg13g2_inv_1 _5707_ (.Y(_2405_),
    .A(_2404_));
 sg13g2_nor2_1 _5708_ (.A(_2400_),
    .B(_2405_),
    .Y(_2406_));
 sg13g2_and2_1 _5709_ (.A(_2400_),
    .B(_2405_),
    .X(_2407_));
 sg13g2_nor3_1 _5710_ (.A(net431),
    .B(net1520),
    .C(_2407_),
    .Y(_0359_));
 sg13g2_a21oi_1 _5711_ (.A1(_2400_),
    .A2(_2405_),
    .Y(_2408_),
    .B1(_2403_));
 sg13g2_a21o_1 _5712_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][11] ),
    .A1(net412),
    .B1(_2401_),
    .X(_2409_));
 sg13g2_nor2b_1 _5713_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][12] ),
    .B_N(_2409_),
    .Y(_2410_));
 sg13g2_xnor2_1 _5714_ (.Y(_2411_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][12] ),
    .B(_2409_));
 sg13g2_nand2_1 _5715_ (.Y(_2412_),
    .A(net1449),
    .B(_2411_));
 sg13g2_xnor2_1 _5716_ (.Y(_2413_),
    .A(net1449),
    .B(_2411_));
 sg13g2_o21ai_1 _5717_ (.B1(net476),
    .Y(_2414_),
    .A1(_2408_),
    .A2(_2413_));
 sg13g2_a21oi_1 _5718_ (.A1(_2408_),
    .A2(net1450),
    .Y(_0360_),
    .B1(_2414_));
 sg13g2_o21ai_1 _5719_ (.B1(_2412_),
    .Y(_2415_),
    .A1(_2408_),
    .A2(_2413_));
 sg13g2_a21oi_2 _5720_ (.B1(_2410_),
    .Y(_2416_),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][12] ),
    .A1(net520));
 sg13g2_and2_1 _5721_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[7] ),
    .B(_2416_),
    .X(_2417_));
 sg13g2_xnor2_1 _5722_ (.Y(_2418_),
    .A(net1549),
    .B(_2416_));
 sg13g2_inv_1 _5723_ (.Y(_2419_),
    .A(_2418_));
 sg13g2_nor2_1 _5724_ (.A(_2415_),
    .B(_2419_),
    .Y(_2420_));
 sg13g2_a21oi_1 _5725_ (.A1(_2415_),
    .A2(_2419_),
    .Y(_2421_),
    .B1(net431));
 sg13g2_nor2b_1 _5726_ (.A(_2420_),
    .B_N(_2421_),
    .Y(_0361_));
 sg13g2_a21oi_1 _5727_ (.A1(_2415_),
    .A2(_2419_),
    .Y(_2422_),
    .B1(_2417_));
 sg13g2_xnor2_1 _5728_ (.Y(_2423_),
    .A(net1117),
    .B(_2416_));
 sg13g2_o21ai_1 _5729_ (.B1(net491),
    .Y(_2424_),
    .A1(_2422_),
    .A2(_2423_));
 sg13g2_a21oi_1 _5730_ (.A1(_2422_),
    .A2(net1118),
    .Y(_0362_),
    .B1(_2424_));
 sg13g2_or2_1 _5731_ (.X(_2425_),
    .B(_2422_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[8] ));
 sg13g2_a21oi_1 _5732_ (.A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[7] ),
    .A2(_2415_),
    .Y(_2426_),
    .B1(_2416_));
 sg13g2_a21oi_1 _5733_ (.A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[8] ),
    .A2(_2416_),
    .Y(_2427_),
    .B1(_2426_));
 sg13g2_a21oi_1 _5734_ (.A1(_2425_),
    .A2(_2427_),
    .Y(_2428_),
    .B1(net903));
 sg13g2_and3_1 _5735_ (.X(_2429_),
    .A(net903),
    .B(_2425_),
    .C(_2427_));
 sg13g2_nor3_1 _5736_ (.A(net431),
    .B(net904),
    .C(_2429_),
    .Y(_0363_));
 sg13g2_nor2_1 _5737_ (.A(net809),
    .B(net427),
    .Y(_0364_));
 sg13g2_nor2b_1 _5738_ (.A(net517),
    .B_N(net877),
    .Y(_2430_));
 sg13g2_xnor2_1 _5739_ (.Y(_2431_),
    .A(net517),
    .B(net877));
 sg13g2_o21ai_1 _5740_ (.B1(net468),
    .Y(_2432_),
    .A1(net809),
    .A2(_2431_));
 sg13g2_a21oi_1 _5741_ (.A1(net809),
    .A2(_2431_),
    .Y(_0365_),
    .B1(_2432_));
 sg13g2_a21oi_1 _5742_ (.A1(net809),
    .A2(_2431_),
    .Y(_2433_),
    .B1(_2430_));
 sg13g2_nand2_1 _5743_ (.Y(_2434_),
    .A(net412),
    .B(net1280));
 sg13g2_xor2_1 _5744_ (.B(net1280),
    .A(net517),
    .X(_2435_));
 sg13g2_o21ai_1 _5745_ (.B1(net468),
    .Y(_2436_),
    .A1(_2433_),
    .A2(_2435_));
 sg13g2_a21oi_1 _5746_ (.A1(_2433_),
    .A2(_2435_),
    .Y(_0366_),
    .B1(_2436_));
 sg13g2_o21ai_1 _5747_ (.B1(_2434_),
    .Y(_2437_),
    .A1(_2433_),
    .A2(_2435_));
 sg13g2_nor2b_1 _5748_ (.A(net517),
    .B_N(net1338),
    .Y(_2438_));
 sg13g2_nand2b_1 _5749_ (.Y(_2439_),
    .B(net517),
    .A_N(net1338));
 sg13g2_nor2b_1 _5750_ (.A(_2438_),
    .B_N(_2439_),
    .Y(_2440_));
 sg13g2_o21ai_1 _5751_ (.B1(net472),
    .Y(_2441_),
    .A1(_2437_),
    .A2(_2440_));
 sg13g2_a21oi_1 _5752_ (.A1(_2437_),
    .A2(_2440_),
    .Y(_0367_),
    .B1(_2441_));
 sg13g2_nand2_1 _5753_ (.Y(_2442_),
    .A(net517),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][4] ));
 sg13g2_xnor2_1 _5754_ (.Y(_2443_),
    .A(net517),
    .B(net1204));
 sg13g2_o21ai_1 _5755_ (.B1(_2439_),
    .Y(_2444_),
    .A1(_2437_),
    .A2(_2438_));
 sg13g2_o21ai_1 _5756_ (.B1(net472),
    .Y(_2445_),
    .A1(_2443_),
    .A2(_2444_));
 sg13g2_a21oi_1 _5757_ (.A1(_2443_),
    .A2(_2444_),
    .Y(_0368_),
    .B1(_2445_));
 sg13g2_o21ai_1 _5758_ (.B1(_2442_),
    .Y(_2446_),
    .A1(_2443_),
    .A2(_2444_));
 sg13g2_nand2b_1 _5759_ (.Y(_2447_),
    .B(net518),
    .A_N(net1084));
 sg13g2_nor2b_1 _5760_ (.A(net517),
    .B_N(net1084),
    .Y(_2448_));
 sg13g2_xnor2_1 _5761_ (.Y(_2449_),
    .A(net518),
    .B(net1084));
 sg13g2_o21ai_1 _5762_ (.B1(net472),
    .Y(_2450_),
    .A1(_2446_),
    .A2(_2449_));
 sg13g2_a21oi_1 _5763_ (.A1(_2446_),
    .A2(_2449_),
    .Y(_0369_),
    .B1(_2450_));
 sg13g2_xnor2_1 _5764_ (.Y(_2451_),
    .A(net518),
    .B(net1354));
 sg13g2_a21oi_1 _5765_ (.A1(_2446_),
    .A2(_2447_),
    .Y(_2452_),
    .B1(_2448_));
 sg13g2_nor2_1 _5766_ (.A(_2451_),
    .B(_2452_),
    .Y(_2453_));
 sg13g2_a21oi_1 _5767_ (.A1(_2451_),
    .A2(_2452_),
    .Y(_2454_),
    .B1(net427));
 sg13g2_nor2b_1 _5768_ (.A(_2453_),
    .B_N(_2454_),
    .Y(_0370_));
 sg13g2_a21oi_1 _5769_ (.A1(net519),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][6] ),
    .Y(_2455_),
    .B1(_2453_));
 sg13g2_nand2_1 _5770_ (.Y(_2456_),
    .A(net412),
    .B(net1078));
 sg13g2_xor2_1 _5771_ (.B(net1078),
    .A(net518),
    .X(_2457_));
 sg13g2_or2_1 _5772_ (.X(_2458_),
    .B(_2457_),
    .A(_2455_));
 sg13g2_nand2_1 _5773_ (.Y(_2459_),
    .A(net461),
    .B(_2458_));
 sg13g2_a21oi_1 _5774_ (.A1(_2455_),
    .A2(_2457_),
    .Y(_0371_),
    .B1(_2459_));
 sg13g2_and2_1 _5775_ (.A(_2456_),
    .B(_2458_),
    .X(_2460_));
 sg13g2_nor2b_1 _5776_ (.A(net519),
    .B_N(net1487),
    .Y(_2461_));
 sg13g2_xor2_1 _5777_ (.B(net1487),
    .A(net519),
    .X(_2462_));
 sg13g2_nor2_1 _5778_ (.A(_2460_),
    .B(_2462_),
    .Y(_2463_));
 sg13g2_a21oi_1 _5779_ (.A1(_2460_),
    .A2(_2462_),
    .Y(_2464_),
    .B1(net425));
 sg13g2_nor2b_1 _5780_ (.A(_2463_),
    .B_N(_2464_),
    .Y(_0372_));
 sg13g2_xnor2_1 _5781_ (.Y(_2465_),
    .A(net520),
    .B(net1127));
 sg13g2_o21ai_1 _5782_ (.B1(_2465_),
    .Y(_2466_),
    .A1(_2461_),
    .A2(_2463_));
 sg13g2_nor3_1 _5783_ (.A(_2461_),
    .B(_2463_),
    .C(_2465_),
    .Y(_2467_));
 sg13g2_nand2_1 _5784_ (.Y(_2468_),
    .A(net476),
    .B(_2466_));
 sg13g2_nor2_1 _5785_ (.A(_2467_),
    .B(_2468_),
    .Y(_0373_));
 sg13g2_a21o_1 _5786_ (.A2(_2465_),
    .A1(_2463_),
    .B1(_2461_),
    .X(_2469_));
 sg13g2_a21oi_1 _5787_ (.A1(_0592_),
    .A2(net1127),
    .Y(_2470_),
    .B1(_2469_));
 sg13g2_xor2_1 _5788_ (.B(net826),
    .A(net520),
    .X(_2471_));
 sg13g2_o21ai_1 _5789_ (.B1(net476),
    .Y(_2472_),
    .A1(_2470_),
    .A2(_2471_));
 sg13g2_a21oi_1 _5790_ (.A1(net1128),
    .A2(_2471_),
    .Y(_0374_),
    .B1(_2472_));
 sg13g2_a21oi_1 _5791_ (.A1(_0592_),
    .A2(net826),
    .Y(_0375_),
    .B1(_2472_));
 sg13g2_and2_1 _5792_ (.A(net1014),
    .B(net1242),
    .X(_2473_));
 sg13g2_o21ai_1 _5793_ (.B1(net457),
    .Y(_2474_),
    .A1(net1014),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[0] ));
 sg13g2_nor2_1 _5794_ (.A(_2473_),
    .B(net1015),
    .Y(_0376_));
 sg13g2_nor2b_1 _5795_ (.A(net512),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[0] ),
    .Y(_2475_));
 sg13g2_xnor2_1 _5796_ (.Y(_2476_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[1] ),
    .B(_2475_));
 sg13g2_nor2_1 _5797_ (.A(_0574_),
    .B(_2476_),
    .Y(_2477_));
 sg13g2_nand2_1 _5798_ (.Y(_2478_),
    .A(_0574_),
    .B(_2476_));
 sg13g2_nor2b_1 _5799_ (.A(_2477_),
    .B_N(_2478_),
    .Y(_2479_));
 sg13g2_nor2_1 _5800_ (.A(_2473_),
    .B(_2479_),
    .Y(_2480_));
 sg13g2_a21oi_1 _5801_ (.A1(_2473_),
    .A2(_2479_),
    .Y(_2481_),
    .B1(net424));
 sg13g2_nor2b_1 _5802_ (.A(net1243),
    .B_N(_2481_),
    .Y(_0377_));
 sg13g2_a21oi_1 _5803_ (.A1(_2473_),
    .A2(_2478_),
    .Y(_2482_),
    .B1(net1428));
 sg13g2_o21ai_1 _5804_ (.B1(net413),
    .Y(_2483_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[0] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[1] ));
 sg13g2_xnor2_1 _5805_ (.Y(_2484_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[2] ),
    .B(_2483_));
 sg13g2_nand2_1 _5806_ (.Y(_2485_),
    .A(net1474),
    .B(_2484_));
 sg13g2_xnor2_1 _5807_ (.Y(_2486_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][2] ),
    .B(_2484_));
 sg13g2_o21ai_1 _5808_ (.B1(net457),
    .Y(_2487_),
    .A1(_2482_),
    .A2(_2486_));
 sg13g2_a21oi_1 _5809_ (.A1(_2482_),
    .A2(_2486_),
    .Y(_0378_),
    .B1(_2487_));
 sg13g2_o21ai_1 _5810_ (.B1(net1475),
    .Y(_2488_),
    .A1(_2482_),
    .A2(_2486_));
 sg13g2_o21ai_1 _5811_ (.B1(_2483_),
    .Y(_2489_),
    .A1(net512),
    .A2(_0575_));
 sg13g2_xor2_1 _5812_ (.B(_2489_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[3] ),
    .X(_2490_));
 sg13g2_and2_1 _5813_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][3] ),
    .B(_2490_),
    .X(_2491_));
 sg13g2_or2_1 _5814_ (.X(_2492_),
    .B(_2490_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][3] ));
 sg13g2_nor2b_1 _5815_ (.A(_2491_),
    .B_N(_2492_),
    .Y(_2493_));
 sg13g2_o21ai_1 _5816_ (.B1(net457),
    .Y(_2494_),
    .A1(_2488_),
    .A2(_2493_));
 sg13g2_a21oi_1 _5817_ (.A1(_2488_),
    .A2(_2493_),
    .Y(_0379_),
    .B1(_2494_));
 sg13g2_a21oi_1 _5818_ (.A1(_2488_),
    .A2(_2492_),
    .Y(_2495_),
    .B1(_2491_));
 sg13g2_nor2b_1 _5819_ (.A(net512),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[3] ),
    .Y(_2496_));
 sg13g2_nor3_1 _5820_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[4] ),
    .B(_2489_),
    .C(_2496_),
    .Y(_2497_));
 sg13g2_o21ai_1 _5821_ (.B1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[4] ),
    .Y(_2498_),
    .A1(_2489_),
    .A2(_2496_));
 sg13g2_nor2b_1 _5822_ (.A(_2497_),
    .B_N(_2498_),
    .Y(_2499_));
 sg13g2_nand2_1 _5823_ (.Y(_2500_),
    .A(net1348),
    .B(_2499_));
 sg13g2_xnor2_1 _5824_ (.Y(_2501_),
    .A(net1348),
    .B(_2499_));
 sg13g2_o21ai_1 _5825_ (.B1(net457),
    .Y(_2502_),
    .A1(_2495_),
    .A2(_2501_));
 sg13g2_a21oi_1 _5826_ (.A1(_2495_),
    .A2(_2501_),
    .Y(_0380_),
    .B1(_2502_));
 sg13g2_o21ai_1 _5827_ (.B1(_2500_),
    .Y(_2503_),
    .A1(_2495_),
    .A2(_2501_));
 sg13g2_nor2_1 _5828_ (.A(net514),
    .B(_2497_),
    .Y(_2504_));
 sg13g2_xnor2_1 _5829_ (.Y(_2505_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[5] ),
    .B(_2504_));
 sg13g2_nor2_1 _5830_ (.A(_0578_),
    .B(_2505_),
    .Y(_2506_));
 sg13g2_nand2_1 _5831_ (.Y(_2507_),
    .A(_0578_),
    .B(_2505_));
 sg13g2_nand2b_1 _5832_ (.Y(_2508_),
    .B(_2507_),
    .A_N(_2506_));
 sg13g2_nor2b_1 _5833_ (.A(_2503_),
    .B_N(_2508_),
    .Y(_2509_));
 sg13g2_nor2b_1 _5834_ (.A(_2508_),
    .B_N(_2503_),
    .Y(_2510_));
 sg13g2_nor3_1 _5835_ (.A(net425),
    .B(_2509_),
    .C(_2510_),
    .Y(_0381_));
 sg13g2_a21oi_1 _5836_ (.A1(_2503_),
    .A2(_2507_),
    .Y(_2511_),
    .B1(_2506_));
 sg13g2_a21o_1 _5837_ (.A2(_2507_),
    .A1(_2503_),
    .B1(_2506_),
    .X(_2512_));
 sg13g2_a21oi_1 _5838_ (.A1(_0577_),
    .A2(_2497_),
    .Y(_2513_),
    .B1(net514));
 sg13g2_xor2_1 _5839_ (.B(_2513_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[6] ),
    .X(_2514_));
 sg13g2_and2_1 _5840_ (.A(net1306),
    .B(_2514_),
    .X(_2515_));
 sg13g2_xnor2_1 _5841_ (.Y(_2516_),
    .A(net1306),
    .B(_2514_));
 sg13g2_inv_1 _5842_ (.Y(_2517_),
    .A(_2516_));
 sg13g2_o21ai_1 _5843_ (.B1(net457),
    .Y(_2518_),
    .A1(_2511_),
    .A2(_2516_));
 sg13g2_a21oi_1 _5844_ (.A1(_2511_),
    .A2(net1307),
    .Y(_0382_),
    .B1(_2518_));
 sg13g2_a21oi_1 _5845_ (.A1(_2512_),
    .A2(_2517_),
    .Y(_2519_),
    .B1(_2515_));
 sg13g2_a21o_1 _5846_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[6] ),
    .A1(net413),
    .B1(_2513_),
    .X(_2520_));
 sg13g2_xor2_1 _5847_ (.B(_2520_),
    .A(net1571),
    .X(_2521_));
 sg13g2_nand2_1 _5848_ (.Y(_2522_),
    .A(net1346),
    .B(_2521_));
 sg13g2_xnor2_1 _5849_ (.Y(_2523_),
    .A(net1346),
    .B(_2521_));
 sg13g2_o21ai_1 _5850_ (.B1(net458),
    .Y(_2524_),
    .A1(_2519_),
    .A2(_2523_));
 sg13g2_a21oi_1 _5851_ (.A1(_2519_),
    .A2(net1347),
    .Y(_0383_),
    .B1(_2524_));
 sg13g2_o21ai_1 _5852_ (.B1(_2522_),
    .Y(_2525_),
    .A1(_2519_),
    .A2(_2523_));
 sg13g2_a21o_1 _5853_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[7] ),
    .A1(net413),
    .B1(_2520_),
    .X(_2526_));
 sg13g2_xnor2_1 _5854_ (.Y(_2527_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[8] ),
    .B(_2526_));
 sg13g2_nor2_1 _5855_ (.A(_0580_),
    .B(_2527_),
    .Y(_2528_));
 sg13g2_nand2_1 _5856_ (.Y(_2529_),
    .A(_0580_),
    .B(_2527_));
 sg13g2_nand2b_1 _5857_ (.Y(_2530_),
    .B(_2529_),
    .A_N(_2528_));
 sg13g2_nand2b_1 _5858_ (.Y(_2531_),
    .B(_2530_),
    .A_N(_2525_));
 sg13g2_nand2b_1 _5859_ (.Y(_2532_),
    .B(_2525_),
    .A_N(_2530_));
 sg13g2_and3_1 _5860_ (.X(_0384_),
    .A(net458),
    .B(_2531_),
    .C(_2532_));
 sg13g2_a21o_1 _5861_ (.A2(_2529_),
    .A1(_2525_),
    .B1(_2528_),
    .X(_2533_));
 sg13g2_a21o_1 _5862_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[8] ),
    .A1(net413),
    .B1(_2526_),
    .X(_2534_));
 sg13g2_xnor2_1 _5863_ (.Y(_2535_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[9] ),
    .B(_2534_));
 sg13g2_nor2b_1 _5864_ (.A(_2535_),
    .B_N(net1326),
    .Y(_2536_));
 sg13g2_xnor2_1 _5865_ (.Y(_2537_),
    .A(net1326),
    .B(_2535_));
 sg13g2_o21ai_1 _5866_ (.B1(net459),
    .Y(_2538_),
    .A1(_2533_),
    .A2(_2537_));
 sg13g2_a21oi_1 _5867_ (.A1(_2533_),
    .A2(net1327),
    .Y(_0385_),
    .B1(_2538_));
 sg13g2_a21oi_1 _5868_ (.A1(_2533_),
    .A2(_2537_),
    .Y(_2539_),
    .B1(_2536_));
 sg13g2_a21oi_1 _5869_ (.A1(net413),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[9] ),
    .Y(_2540_),
    .B1(_2534_));
 sg13g2_xnor2_1 _5870_ (.Y(_2541_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[10] ),
    .B(_2540_));
 sg13g2_nand2_1 _5871_ (.Y(_2542_),
    .A(net1422),
    .B(_2541_));
 sg13g2_xnor2_1 _5872_ (.Y(_2543_),
    .A(net1422),
    .B(_2541_));
 sg13g2_o21ai_1 _5873_ (.B1(net459),
    .Y(_2544_),
    .A1(_2539_),
    .A2(_2543_));
 sg13g2_a21oi_1 _5874_ (.A1(_2539_),
    .A2(net1423),
    .Y(_0386_),
    .B1(_2544_));
 sg13g2_o21ai_1 _5875_ (.B1(_2542_),
    .Y(_2545_),
    .A1(_2539_),
    .A2(_2543_));
 sg13g2_nand2_1 _5876_ (.Y(_2546_),
    .A(net513),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[10] ));
 sg13g2_o21ai_1 _5877_ (.B1(_2546_),
    .Y(_2547_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[10] ),
    .A2(_2540_));
 sg13g2_and2_1 _5878_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][11] ),
    .B(_2547_),
    .X(_2548_));
 sg13g2_xor2_1 _5879_ (.B(_2547_),
    .A(net1486),
    .X(_2549_));
 sg13g2_o21ai_1 _5880_ (.B1(net459),
    .Y(_2550_),
    .A1(_2545_),
    .A2(_2549_));
 sg13g2_a21oi_1 _5881_ (.A1(_2545_),
    .A2(_2549_),
    .Y(_0387_),
    .B1(_2550_));
 sg13g2_a21oi_1 _5882_ (.A1(_2545_),
    .A2(_2549_),
    .Y(_2551_),
    .B1(_2548_));
 sg13g2_xnor2_1 _5883_ (.Y(_2552_),
    .A(net1217),
    .B(_2547_));
 sg13g2_o21ai_1 _5884_ (.B1(net459),
    .Y(_2553_),
    .A1(_2551_),
    .A2(_2552_));
 sg13g2_a21oi_1 _5885_ (.A1(_2551_),
    .A2(_2552_),
    .Y(_0388_),
    .B1(_2553_));
 sg13g2_nor2b_1 _5886_ (.A(net973),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][2] ),
    .Y(_2554_));
 sg13g2_xnor2_1 _5887_ (.Y(_2555_),
    .A(net973),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][2] ));
 sg13g2_nor2_1 _5888_ (.A(net425),
    .B(net974),
    .Y(_0389_));
 sg13g2_nor2b_1 _5889_ (.A(net512),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][2] ),
    .Y(_2556_));
 sg13g2_xnor2_1 _5890_ (.Y(_2557_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][3] ),
    .B(_2556_));
 sg13g2_nand2_1 _5891_ (.Y(_2558_),
    .A(net1146),
    .B(_2557_));
 sg13g2_xnor2_1 _5892_ (.Y(_2559_),
    .A(net1146),
    .B(_2557_));
 sg13g2_o21ai_1 _5893_ (.B1(net457),
    .Y(_2560_),
    .A1(_2554_),
    .A2(_2559_));
 sg13g2_a21oi_1 _5894_ (.A1(_2554_),
    .A2(net1147),
    .Y(_0390_),
    .B1(_2560_));
 sg13g2_o21ai_1 _5895_ (.B1(_2558_),
    .Y(_2561_),
    .A1(_2554_),
    .A2(_2559_));
 sg13g2_o21ai_1 _5896_ (.B1(net413),
    .Y(_2562_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][2] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][3] ));
 sg13g2_xnor2_1 _5897_ (.Y(_2563_),
    .A(net1481),
    .B(_2562_));
 sg13g2_nor2b_1 _5898_ (.A(_2563_),
    .B_N(net1242),
    .Y(_2564_));
 sg13g2_xnor2_1 _5899_ (.Y(_2565_),
    .A(net1242),
    .B(_2563_));
 sg13g2_nor2_1 _5900_ (.A(_2561_),
    .B(_2565_),
    .Y(_2566_));
 sg13g2_a21oi_1 _5901_ (.A1(_2561_),
    .A2(_2565_),
    .Y(_2567_),
    .B1(net424));
 sg13g2_nor2b_1 _5902_ (.A(_2566_),
    .B_N(_2567_),
    .Y(_0391_));
 sg13g2_a21o_1 _5903_ (.A2(_2565_),
    .A1(_2561_),
    .B1(_2564_),
    .X(_2568_));
 sg13g2_o21ai_1 _5904_ (.B1(_2562_),
    .Y(_2569_),
    .A1(net512),
    .A2(_0576_));
 sg13g2_xnor2_1 _5905_ (.Y(_2570_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][5] ),
    .B(_2569_));
 sg13g2_and2_1 _5906_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[1] ),
    .B(_2570_),
    .X(_2571_));
 sg13g2_xor2_1 _5907_ (.B(_2570_),
    .A(net1509),
    .X(_2572_));
 sg13g2_o21ai_1 _5908_ (.B1(net457),
    .Y(_2573_),
    .A1(_2568_),
    .A2(_2572_));
 sg13g2_a21oi_1 _5909_ (.A1(_2568_),
    .A2(net1510),
    .Y(_0392_),
    .B1(_2573_));
 sg13g2_a21oi_1 _5910_ (.A1(_2568_),
    .A2(_2572_),
    .Y(_2574_),
    .B1(_2571_));
 sg13g2_and3_1 _5911_ (.X(_2575_),
    .A(_0576_),
    .B(_0578_),
    .C(_2562_));
 sg13g2_nor2_1 _5912_ (.A(net512),
    .B(_2575_),
    .Y(_2576_));
 sg13g2_xnor2_1 _5913_ (.Y(_2577_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][6] ),
    .B(_2576_));
 sg13g2_nand2_1 _5914_ (.Y(_2578_),
    .A(net1248),
    .B(_2577_));
 sg13g2_nor2_1 _5915_ (.A(net1248),
    .B(_2577_),
    .Y(_2579_));
 sg13g2_xnor2_1 _5916_ (.Y(_2580_),
    .A(net1248),
    .B(_2577_));
 sg13g2_o21ai_1 _5917_ (.B1(net457),
    .Y(_2581_),
    .A1(_2574_),
    .A2(_2580_));
 sg13g2_a21oi_1 _5918_ (.A1(_2574_),
    .A2(net1249),
    .Y(_0393_),
    .B1(_2581_));
 sg13g2_o21ai_1 _5919_ (.B1(_2578_),
    .Y(_2582_),
    .A1(_2574_),
    .A2(_2579_));
 sg13g2_a21oi_1 _5920_ (.A1(_0579_),
    .A2(_2575_),
    .Y(_2583_),
    .B1(net512));
 sg13g2_xnor2_1 _5921_ (.Y(_2584_),
    .A(net1346),
    .B(_2583_));
 sg13g2_and2_1 _5922_ (.A(net1381),
    .B(_2584_),
    .X(_2585_));
 sg13g2_xnor2_1 _5923_ (.Y(_2586_),
    .A(net1381),
    .B(_2584_));
 sg13g2_inv_1 _5924_ (.Y(_2587_),
    .A(_2586_));
 sg13g2_o21ai_1 _5925_ (.B1(net458),
    .Y(_2588_),
    .A1(_2582_),
    .A2(_2587_));
 sg13g2_a21oi_1 _5926_ (.A1(_2582_),
    .A2(_2587_),
    .Y(_0394_),
    .B1(_2588_));
 sg13g2_a21o_1 _5927_ (.A2(_2587_),
    .A1(_2582_),
    .B1(_2585_),
    .X(_2589_));
 sg13g2_a21oi_1 _5928_ (.A1(net413),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][7] ),
    .Y(_2590_),
    .B1(_2583_));
 sg13g2_xnor2_1 _5929_ (.Y(_2591_),
    .A(net1575),
    .B(_2590_));
 sg13g2_nor2b_1 _5930_ (.A(_2591_),
    .B_N(net1454),
    .Y(_2592_));
 sg13g2_xnor2_1 _5931_ (.Y(_2593_),
    .A(net1454),
    .B(_2591_));
 sg13g2_nor2_1 _5932_ (.A(_2589_),
    .B(net1455),
    .Y(_2594_));
 sg13g2_and2_1 _5933_ (.A(_2589_),
    .B(_2593_),
    .X(_2595_));
 sg13g2_nor3_1 _5934_ (.A(net425),
    .B(_2594_),
    .C(_2595_),
    .Y(_0395_));
 sg13g2_a21o_1 _5935_ (.A2(_2593_),
    .A1(_2589_),
    .B1(_2592_),
    .X(_2596_));
 sg13g2_o21ai_1 _5936_ (.B1(_2590_),
    .Y(_2597_),
    .A1(net514),
    .A2(_0580_));
 sg13g2_xnor2_1 _5937_ (.Y(_2598_),
    .A(net1326),
    .B(_2597_));
 sg13g2_and2_1 _5938_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[5] ),
    .B(_2598_),
    .X(_2599_));
 sg13g2_xnor2_1 _5939_ (.Y(_2600_),
    .A(_0577_),
    .B(_2598_));
 sg13g2_o21ai_1 _5940_ (.B1(net458),
    .Y(_2601_),
    .A1(_2596_),
    .A2(_2600_));
 sg13g2_a21oi_1 _5941_ (.A1(_2596_),
    .A2(_2600_),
    .Y(_0396_),
    .B1(_2601_));
 sg13g2_a21oi_1 _5942_ (.A1(_2596_),
    .A2(_2600_),
    .Y(_2602_),
    .B1(_2599_));
 sg13g2_a21o_1 _5943_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][9] ),
    .A1(net413),
    .B1(_2597_),
    .X(_2603_));
 sg13g2_xnor2_1 _5944_ (.Y(_2604_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][10] ),
    .B(_2603_));
 sg13g2_nand2_1 _5945_ (.Y(_2605_),
    .A(net1435),
    .B(_2604_));
 sg13g2_xnor2_1 _5946_ (.Y(_2606_),
    .A(net1435),
    .B(_2604_));
 sg13g2_o21ai_1 _5947_ (.B1(net459),
    .Y(_2607_),
    .A1(_2602_),
    .A2(_2606_));
 sg13g2_a21oi_1 _5948_ (.A1(_2602_),
    .A2(net1436),
    .Y(_0397_),
    .B1(_2607_));
 sg13g2_o21ai_1 _5949_ (.B1(_2605_),
    .Y(_2608_),
    .A1(_2602_),
    .A2(_2606_));
 sg13g2_a21o_1 _5950_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][10] ),
    .A1(net414),
    .B1(_2603_),
    .X(_2609_));
 sg13g2_xnor2_1 _5951_ (.Y(_2610_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][11] ),
    .B(_2609_));
 sg13g2_nand2_1 _5952_ (.Y(_2611_),
    .A(net1457),
    .B(_2610_));
 sg13g2_xor2_1 _5953_ (.B(_2610_),
    .A(net1457),
    .X(_2612_));
 sg13g2_nand2_1 _5954_ (.Y(_2613_),
    .A(_2608_),
    .B(_2612_));
 sg13g2_o21ai_1 _5955_ (.B1(net459),
    .Y(_2614_),
    .A1(_2608_),
    .A2(_2612_));
 sg13g2_nor2b_1 _5956_ (.A(_2614_),
    .B_N(_2613_),
    .Y(_0398_));
 sg13g2_a21o_1 _5957_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][11] ),
    .A1(net414),
    .B1(_2609_),
    .X(_2615_));
 sg13g2_xnor2_1 _5958_ (.Y(_2616_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][12] ),
    .B(_2615_));
 sg13g2_nand2_1 _5959_ (.Y(_2617_),
    .A(net1530),
    .B(_2616_));
 sg13g2_xnor2_1 _5960_ (.Y(_2618_),
    .A(net1530),
    .B(_2616_));
 sg13g2_and3_1 _5961_ (.X(_2619_),
    .A(_2611_),
    .B(_2613_),
    .C(_2618_));
 sg13g2_a21oi_1 _5962_ (.A1(_2611_),
    .A2(_2613_),
    .Y(_2620_),
    .B1(_2618_));
 sg13g2_a21o_1 _5963_ (.A2(_2613_),
    .A1(_2611_),
    .B1(_2618_),
    .X(_2621_));
 sg13g2_nor3_1 _5964_ (.A(net425),
    .B(_2619_),
    .C(_2620_),
    .Y(_0399_));
 sg13g2_mux2_1 _5965_ (.A0(_2615_),
    .A1(net513),
    .S(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][12] ),
    .X(_2622_));
 sg13g2_nand2_1 _5966_ (.Y(_2623_),
    .A(_0581_),
    .B(_2622_));
 sg13g2_xnor2_1 _5967_ (.Y(_2624_),
    .A(_0581_),
    .B(_2622_));
 sg13g2_and3_1 _5968_ (.X(_2625_),
    .A(_2617_),
    .B(_2621_),
    .C(_2624_));
 sg13g2_a21oi_1 _5969_ (.A1(_2617_),
    .A2(_2621_),
    .Y(_2626_),
    .B1(_2624_));
 sg13g2_nor3_1 _5970_ (.A(net425),
    .B(_2625_),
    .C(_2626_),
    .Y(_0400_));
 sg13g2_o21ai_1 _5971_ (.B1(_2617_),
    .Y(_2627_),
    .A1(_0581_),
    .A2(_2622_));
 sg13g2_a21oi_1 _5972_ (.A1(_2620_),
    .A2(_2623_),
    .Y(_2628_),
    .B1(_2627_));
 sg13g2_xor2_1 _5973_ (.B(_2622_),
    .A(net1323),
    .X(_2629_));
 sg13g2_o21ai_1 _5974_ (.B1(net459),
    .Y(_2630_),
    .A1(_2628_),
    .A2(_2629_));
 sg13g2_a21oi_1 _5975_ (.A1(_2628_),
    .A2(_2629_),
    .Y(_0401_),
    .B1(_2630_));
 sg13g2_and2_1 _5976_ (.A(net467),
    .B(net791),
    .X(_0402_));
 sg13g2_and2_1 _5977_ (.A(net467),
    .B(net768),
    .X(_0403_));
 sg13g2_and2_1 _5978_ (.A(net467),
    .B(net766),
    .X(_0404_));
 sg13g2_and2_1 _5979_ (.A(net467),
    .B(net783),
    .X(_0405_));
 sg13g2_and2_1 _5980_ (.A(net467),
    .B(net773),
    .X(_0406_));
 sg13g2_nor2_1 _5981_ (.A(net810),
    .B(net427),
    .Y(_0407_));
 sg13g2_nor2b_1 _5982_ (.A(net513),
    .B_N(net841),
    .Y(_2631_));
 sg13g2_xnor2_1 _5983_ (.Y(_2632_),
    .A(net513),
    .B(net841));
 sg13g2_o21ai_1 _5984_ (.B1(net467),
    .Y(_2633_),
    .A1(net810),
    .A2(_2632_));
 sg13g2_a21oi_1 _5985_ (.A1(net810),
    .A2(_2632_),
    .Y(_0408_),
    .B1(_2633_));
 sg13g2_a21oi_1 _5986_ (.A1(net810),
    .A2(_2632_),
    .Y(_2634_),
    .B1(_2631_));
 sg13g2_nand2_1 _5987_ (.Y(_2635_),
    .A(net513),
    .B(net1051));
 sg13g2_xnor2_1 _5988_ (.Y(_2636_),
    .A(net513),
    .B(net1051));
 sg13g2_or2_1 _5989_ (.X(_2637_),
    .B(_2636_),
    .A(_2634_));
 sg13g2_nand2_1 _5990_ (.Y(_2638_),
    .A(net460),
    .B(_2637_));
 sg13g2_a21oi_1 _5991_ (.A1(_2634_),
    .A2(_2636_),
    .Y(_0409_),
    .B1(_2638_));
 sg13g2_nand2_1 _5992_ (.Y(_2639_),
    .A(net414),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][8] ));
 sg13g2_xor2_1 _5993_ (.B(net1325),
    .A(net513),
    .X(_2640_));
 sg13g2_nand3_1 _5994_ (.B(_2637_),
    .C(_2640_),
    .A(_2635_),
    .Y(_2641_));
 sg13g2_a21o_1 _5995_ (.A2(_2637_),
    .A1(_2635_),
    .B1(_2640_),
    .X(_2642_));
 sg13g2_and3_1 _5996_ (.X(_0410_),
    .A(net460),
    .B(_2641_),
    .C(_2642_));
 sg13g2_and2_1 _5997_ (.A(_2639_),
    .B(_2642_),
    .X(_2643_));
 sg13g2_xor2_1 _5998_ (.B(net1154),
    .A(net513),
    .X(_2644_));
 sg13g2_or2_1 _5999_ (.X(_2645_),
    .B(_2644_),
    .A(_2643_));
 sg13g2_nand2_1 _6000_ (.Y(_2646_),
    .A(net460),
    .B(_2645_));
 sg13g2_a21oi_1 _6001_ (.A1(_2643_),
    .A2(_2644_),
    .Y(_0411_),
    .B1(_2646_));
 sg13g2_o21ai_1 _6002_ (.B1(_2645_),
    .Y(_2647_),
    .A1(net514),
    .A2(_0588_));
 sg13g2_xnor2_1 _6003_ (.Y(_2648_),
    .A(net514),
    .B(net1068));
 sg13g2_o21ai_1 _6004_ (.B1(net460),
    .Y(_2649_),
    .A1(_2647_),
    .A2(_2648_));
 sg13g2_a21oi_1 _6005_ (.A1(_2647_),
    .A2(_2648_),
    .Y(_0412_),
    .B1(_2649_));
 sg13g2_nand2b_1 _6006_ (.Y(_2650_),
    .B(_2648_),
    .A_N(_2645_));
 sg13g2_o21ai_1 _6007_ (.B1(net414),
    .Y(_2651_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][9] ),
    .A2(net1068));
 sg13g2_and3_1 _6008_ (.X(_0413_),
    .A(net460),
    .B(_2650_),
    .C(net1069));
 sg13g2_nand2_1 _6009_ (.Y(_2652_),
    .A(net1046),
    .B(net1076));
 sg13g2_o21ai_1 _6010_ (.B1(net452),
    .Y(_2653_),
    .A1(net1046),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[0] ));
 sg13g2_nor2b_1 _6011_ (.A(net1047),
    .B_N(_2652_),
    .Y(_0414_));
 sg13g2_nor2b_1 _6012_ (.A(net507),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[0] ),
    .Y(_2654_));
 sg13g2_xnor2_1 _6013_ (.Y(_2655_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[1] ),
    .B(_2654_));
 sg13g2_or2_1 _6014_ (.X(_2656_),
    .B(_2655_),
    .A(_0545_));
 sg13g2_xnor2_1 _6015_ (.Y(_2657_),
    .A(_0545_),
    .B(_2655_));
 sg13g2_o21ai_1 _6016_ (.B1(net452),
    .Y(_2658_),
    .A1(_2652_),
    .A2(_2657_));
 sg13g2_a21oi_1 _6017_ (.A1(_2652_),
    .A2(_2657_),
    .Y(_0415_),
    .B1(_2658_));
 sg13g2_o21ai_1 _6018_ (.B1(_2656_),
    .Y(_2659_),
    .A1(_2652_),
    .A2(_2657_));
 sg13g2_o21ai_1 _6019_ (.B1(net416),
    .Y(_2660_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[0] ),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[1] ));
 sg13g2_xnor2_1 _6020_ (.Y(_2661_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[2] ),
    .B(_2660_));
 sg13g2_and2_1 _6021_ (.A(net1264),
    .B(_2661_),
    .X(_2662_));
 sg13g2_or2_1 _6022_ (.X(_2663_),
    .B(_2661_),
    .A(net1264));
 sg13g2_nor2b_1 _6023_ (.A(_2662_),
    .B_N(_2663_),
    .Y(_2664_));
 sg13g2_nor2_1 _6024_ (.A(_2659_),
    .B(_2664_),
    .Y(_2665_));
 sg13g2_a21oi_1 _6025_ (.A1(_2659_),
    .A2(_2664_),
    .Y(_2666_),
    .B1(net422));
 sg13g2_nor2b_1 _6026_ (.A(_2665_),
    .B_N(_2666_),
    .Y(_0416_));
 sg13g2_a21oi_1 _6027_ (.A1(_2659_),
    .A2(_2663_),
    .Y(_2667_),
    .B1(_2662_));
 sg13g2_nor3_1 _6028_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[0] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[1] ),
    .C(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[2] ),
    .Y(_2668_));
 sg13g2_nor2_1 _6029_ (.A(net507),
    .B(_2668_),
    .Y(_2669_));
 sg13g2_xnor2_1 _6030_ (.Y(_2670_),
    .A(_0620_),
    .B(_2669_));
 sg13g2_nand2_1 _6031_ (.Y(_2671_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][3] ),
    .B(_2670_));
 sg13g2_xnor2_1 _6032_ (.Y(_2672_),
    .A(net1339),
    .B(_2670_));
 sg13g2_or2_1 _6033_ (.X(_2673_),
    .B(_2672_),
    .A(_2667_));
 sg13g2_nand2_1 _6034_ (.Y(_2674_),
    .A(net452),
    .B(_2673_));
 sg13g2_a21oi_1 _6035_ (.A1(_2667_),
    .A2(_2672_),
    .Y(_0417_),
    .B1(_2674_));
 sg13g2_and2_1 _6036_ (.A(_2671_),
    .B(_2673_),
    .X(_2675_));
 sg13g2_o21ai_1 _6037_ (.B1(_2671_),
    .Y(_2676_),
    .A1(_2667_),
    .A2(_2672_));
 sg13g2_a21oi_1 _6038_ (.A1(_0620_),
    .A2(_2668_),
    .Y(_2677_),
    .B1(net507));
 sg13g2_xor2_1 _6039_ (.B(_2677_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[4] ),
    .X(_2678_));
 sg13g2_and2_1 _6040_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][4] ),
    .B(_2678_),
    .X(_2679_));
 sg13g2_xnor2_1 _6041_ (.Y(_2680_),
    .A(net1295),
    .B(_2678_));
 sg13g2_inv_1 _6042_ (.Y(_2681_),
    .A(_2680_));
 sg13g2_o21ai_1 _6043_ (.B1(net452),
    .Y(_2682_),
    .A1(_2675_),
    .A2(_2680_));
 sg13g2_a21oi_1 _6044_ (.A1(_2675_),
    .A2(net1296),
    .Y(_0418_),
    .B1(_2682_));
 sg13g2_a21oi_1 _6045_ (.A1(_2676_),
    .A2(_2681_),
    .Y(_2683_),
    .B1(_2679_));
 sg13g2_a21o_1 _6046_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[4] ),
    .A1(net416),
    .B1(_2677_),
    .X(_2684_));
 sg13g2_xor2_1 _6047_ (.B(_2684_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[5] ),
    .X(_2685_));
 sg13g2_nor2_1 _6048_ (.A(net1209),
    .B(_2685_),
    .Y(_2686_));
 sg13g2_xnor2_1 _6049_ (.Y(_2687_),
    .A(net1209),
    .B(_2685_));
 sg13g2_o21ai_1 _6050_ (.B1(net452),
    .Y(_2688_),
    .A1(_2683_),
    .A2(_2687_));
 sg13g2_a21oi_1 _6051_ (.A1(_2683_),
    .A2(net1210),
    .Y(_0419_),
    .B1(_2688_));
 sg13g2_a21oi_1 _6052_ (.A1(net416),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[5] ),
    .Y(_2689_),
    .B1(_2684_));
 sg13g2_xnor2_1 _6053_ (.Y(_2690_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[6] ),
    .B(_2689_));
 sg13g2_and2_1 _6054_ (.A(net1522),
    .B(_2690_),
    .X(_2691_));
 sg13g2_xnor2_1 _6055_ (.Y(_2692_),
    .A(net1522),
    .B(_2690_));
 sg13g2_a221oi_1 _6056_ (.B2(net1209),
    .C1(_2679_),
    .B1(_2685_),
    .A1(_2676_),
    .Y(_2693_),
    .A2(_2681_));
 sg13g2_o21ai_1 _6057_ (.B1(_2692_),
    .Y(_2694_),
    .A1(_2686_),
    .A2(_2693_));
 sg13g2_nor3_1 _6058_ (.A(_2686_),
    .B(_2692_),
    .C(_2693_),
    .Y(_2695_));
 sg13g2_nor2_1 _6059_ (.A(net424),
    .B(_2695_),
    .Y(_2696_));
 sg13g2_and2_1 _6060_ (.A(net1523),
    .B(_2696_),
    .X(_0420_));
 sg13g2_nand2_1 _6061_ (.Y(_2697_),
    .A(net416),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[6] ));
 sg13g2_and2_1 _6062_ (.A(_2689_),
    .B(_2697_),
    .X(_2698_));
 sg13g2_xnor2_1 _6063_ (.Y(_2699_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[7] ),
    .B(_2698_));
 sg13g2_nand2_1 _6064_ (.Y(_2700_),
    .A(net1318),
    .B(_2699_));
 sg13g2_xnor2_1 _6065_ (.Y(_2701_),
    .A(net1318),
    .B(_2699_));
 sg13g2_inv_1 _6066_ (.Y(_2702_),
    .A(_2701_));
 sg13g2_nor3_1 _6067_ (.A(_2691_),
    .B(_2695_),
    .C(_2702_),
    .Y(_2703_));
 sg13g2_o21ai_1 _6068_ (.B1(_2702_),
    .Y(_2704_),
    .A1(_2691_),
    .A2(_2695_));
 sg13g2_nand2_1 _6069_ (.Y(_2705_),
    .A(net452),
    .B(_2704_));
 sg13g2_nor2_1 _6070_ (.A(_2703_),
    .B(_2705_),
    .Y(_0421_));
 sg13g2_o21ai_1 _6071_ (.B1(_2698_),
    .Y(_2706_),
    .A1(net511),
    .A2(_0622_));
 sg13g2_xnor2_1 _6072_ (.Y(_2707_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[8] ),
    .B(_2706_));
 sg13g2_nand2b_1 _6073_ (.Y(_2708_),
    .B(net1497),
    .A_N(_2707_));
 sg13g2_xor2_1 _6074_ (.B(_2707_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][8] ),
    .X(_2709_));
 sg13g2_nand3_1 _6075_ (.B(_2704_),
    .C(_2709_),
    .A(net1319),
    .Y(_2710_));
 sg13g2_a21o_1 _6076_ (.A2(_2704_),
    .A1(_2700_),
    .B1(_2709_),
    .X(_2711_));
 sg13g2_and3_1 _6077_ (.X(_0422_),
    .A(net453),
    .B(net1320),
    .C(_2711_));
 sg13g2_a21o_1 _6078_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[8] ),
    .A1(net416),
    .B1(_2706_),
    .X(_2712_));
 sg13g2_xnor2_1 _6079_ (.Y(_2713_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[9] ),
    .B(_2712_));
 sg13g2_nand2b_1 _6080_ (.Y(_2714_),
    .B(net1371),
    .A_N(_2713_));
 sg13g2_xnor2_1 _6081_ (.Y(_2715_),
    .A(_0623_),
    .B(_2713_));
 sg13g2_nand3_1 _6082_ (.B(_2711_),
    .C(_2715_),
    .A(_2708_),
    .Y(_2716_));
 sg13g2_a21o_1 _6083_ (.A2(_2711_),
    .A1(_2708_),
    .B1(_2715_),
    .X(_2717_));
 sg13g2_and3_1 _6084_ (.X(_0423_),
    .A(net454),
    .B(net1498),
    .C(_2717_));
 sg13g2_a21oi_1 _6085_ (.A1(net417),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[9] ),
    .Y(_2718_),
    .B1(_2712_));
 sg13g2_xnor2_1 _6086_ (.Y(_2719_),
    .A(_0625_),
    .B(_2718_));
 sg13g2_nor2b_1 _6087_ (.A(_2719_),
    .B_N(net1557),
    .Y(_2720_));
 sg13g2_xor2_1 _6088_ (.B(_2719_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][10] ),
    .X(_2721_));
 sg13g2_and3_1 _6089_ (.X(_2722_),
    .A(_2714_),
    .B(_2717_),
    .C(_2721_));
 sg13g2_a21oi_1 _6090_ (.A1(_2714_),
    .A2(_2717_),
    .Y(_2723_),
    .B1(_2721_));
 sg13g2_nor3_1 _6091_ (.A(net424),
    .B(net1372),
    .C(_2723_),
    .Y(_0424_));
 sg13g2_o21ai_1 _6092_ (.B1(_2718_),
    .Y(_2724_),
    .A1(net510),
    .A2(_0625_));
 sg13g2_xor2_1 _6093_ (.B(_2724_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[11] ),
    .X(_2725_));
 sg13g2_nand2_1 _6094_ (.Y(_2726_),
    .A(net1130),
    .B(_2725_));
 sg13g2_xnor2_1 _6095_ (.Y(_2727_),
    .A(_0624_),
    .B(_2725_));
 sg13g2_nor3_1 _6096_ (.A(_2720_),
    .B(_2723_),
    .C(_2727_),
    .Y(_2728_));
 sg13g2_o21ai_1 _6097_ (.B1(_2727_),
    .Y(_2729_),
    .A1(_2720_),
    .A2(_2723_));
 sg13g2_nand2_1 _6098_ (.Y(_2730_),
    .A(net454),
    .B(_2729_));
 sg13g2_nor2_1 _6099_ (.A(_2728_),
    .B(_2730_),
    .Y(_0425_));
 sg13g2_nand2_1 _6100_ (.Y(_2731_),
    .A(net1131),
    .B(_2729_));
 sg13g2_mux2_1 _6101_ (.A0(_2724_),
    .A1(net510),
    .S(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[11] ),
    .X(_2732_));
 sg13g2_xor2_1 _6102_ (.B(_2732_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][12] ),
    .X(_2733_));
 sg13g2_o21ai_1 _6103_ (.B1(net454),
    .Y(_2734_),
    .A1(_2731_),
    .A2(_2733_));
 sg13g2_a21oi_1 _6104_ (.A1(_2731_),
    .A2(_2733_),
    .Y(_0426_),
    .B1(_2734_));
 sg13g2_nor2_1 _6105_ (.A(net1046),
    .B(_0545_),
    .Y(_2735_));
 sg13g2_xnor2_1 _6106_ (.Y(_2736_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][0] ),
    .B(net965));
 sg13g2_nor2_1 _6107_ (.A(net424),
    .B(net966),
    .Y(_0427_));
 sg13g2_nor2b_1 _6108_ (.A(net507),
    .B_N(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][1] ),
    .Y(_2737_));
 sg13g2_xnor2_1 _6109_ (.Y(_2738_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][2] ),
    .B(_2737_));
 sg13g2_nand2_1 _6110_ (.Y(_2739_),
    .A(net1076),
    .B(_2738_));
 sg13g2_xnor2_1 _6111_ (.Y(_2740_),
    .A(net1076),
    .B(net1265));
 sg13g2_o21ai_1 _6112_ (.B1(net452),
    .Y(_2741_),
    .A1(_2735_),
    .A2(_2740_));
 sg13g2_a21oi_1 _6113_ (.A1(_2735_),
    .A2(_2740_),
    .Y(_0428_),
    .B1(_2741_));
 sg13g2_o21ai_1 _6114_ (.B1(_2739_),
    .Y(_2742_),
    .A1(_2735_),
    .A2(_2740_));
 sg13g2_nor2_1 _6115_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][1] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][2] ),
    .Y(_2743_));
 sg13g2_nor2_1 _6116_ (.A(net507),
    .B(_2743_),
    .Y(_2744_));
 sg13g2_xnor2_1 _6117_ (.Y(_2745_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][3] ),
    .B(_2744_));
 sg13g2_and2_1 _6118_ (.A(net1552),
    .B(_2745_),
    .X(_2746_));
 sg13g2_or2_1 _6119_ (.X(_2747_),
    .B(_2745_),
    .A(net1552));
 sg13g2_nor2b_1 _6120_ (.A(_2746_),
    .B_N(_2747_),
    .Y(_2748_));
 sg13g2_nor2_1 _6121_ (.A(_2742_),
    .B(_2748_),
    .Y(_2749_));
 sg13g2_a21oi_1 _6122_ (.A1(_2742_),
    .A2(_2748_),
    .Y(_2750_),
    .B1(net422));
 sg13g2_nor2b_1 _6123_ (.A(_2749_),
    .B_N(_2750_),
    .Y(_0429_));
 sg13g2_a21o_1 _6124_ (.A2(_2747_),
    .A1(_2742_),
    .B1(_2746_),
    .X(_2751_));
 sg13g2_a21oi_1 _6125_ (.A1(_0619_),
    .A2(_2743_),
    .Y(_2752_),
    .B1(net507));
 sg13g2_xor2_1 _6126_ (.B(_2752_),
    .A(net1295),
    .X(_2753_));
 sg13g2_nor2b_1 _6127_ (.A(_2753_),
    .B_N(net1298),
    .Y(_2754_));
 sg13g2_xnor2_1 _6128_ (.Y(_2755_),
    .A(net1298),
    .B(_2753_));
 sg13g2_o21ai_1 _6129_ (.B1(net452),
    .Y(_2756_),
    .A1(_2751_),
    .A2(_2755_));
 sg13g2_a21oi_1 _6130_ (.A1(_2751_),
    .A2(_2755_),
    .Y(_0430_),
    .B1(_2756_));
 sg13g2_a21o_1 _6131_ (.A2(_2755_),
    .A1(_2751_),
    .B1(_2754_),
    .X(_2757_));
 sg13g2_a21o_1 _6132_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][4] ),
    .A1(net416),
    .B1(_2752_),
    .X(_2758_));
 sg13g2_xnor2_1 _6133_ (.Y(_2759_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][5] ),
    .B(_2758_));
 sg13g2_and2_1 _6134_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[3] ),
    .B(_2759_),
    .X(_2760_));
 sg13g2_xnor2_1 _6135_ (.Y(_2761_),
    .A(_0620_),
    .B(_2759_));
 sg13g2_nor2_1 _6136_ (.A(_2757_),
    .B(net1547),
    .Y(_2762_));
 sg13g2_a21oi_1 _6137_ (.A1(_2757_),
    .A2(_2761_),
    .Y(_2763_),
    .B1(net422));
 sg13g2_nor2b_1 _6138_ (.A(_2762_),
    .B_N(_2763_),
    .Y(_0431_));
 sg13g2_a21oi_1 _6139_ (.A1(_2757_),
    .A2(_2761_),
    .Y(_2764_),
    .B1(_2760_));
 sg13g2_a21o_1 _6140_ (.A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][5] ),
    .A1(net416),
    .B1(_2758_),
    .X(_2765_));
 sg13g2_xnor2_1 _6141_ (.Y(_2766_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][6] ),
    .B(_2765_));
 sg13g2_nand2_1 _6142_ (.Y(_2767_),
    .A(net1406),
    .B(_2766_));
 sg13g2_xnor2_1 _6143_ (.Y(_2768_),
    .A(net1406),
    .B(_2766_));
 sg13g2_o21ai_1 _6144_ (.B1(net453),
    .Y(_2769_),
    .A1(_2764_),
    .A2(_2768_));
 sg13g2_a21oi_1 _6145_ (.A1(_2764_),
    .A2(_2768_),
    .Y(_0432_),
    .B1(_2769_));
 sg13g2_o21ai_1 _6146_ (.B1(_2767_),
    .Y(_2770_),
    .A1(_2764_),
    .A2(_2768_));
 sg13g2_inv_1 _6147_ (.Y(_2771_),
    .A(_2770_));
 sg13g2_a21oi_1 _6148_ (.A1(net416),
    .A2(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][6] ),
    .Y(_2772_),
    .B1(_2765_));
 sg13g2_xnor2_1 _6149_ (.Y(_2773_),
    .A(_0621_),
    .B(_2772_));
 sg13g2_and2_1 _6150_ (.A(net1420),
    .B(_2773_),
    .X(_2774_));
 sg13g2_xnor2_1 _6151_ (.Y(_2775_),
    .A(net1420),
    .B(_2773_));
 sg13g2_inv_1 _6152_ (.Y(_2776_),
    .A(_2775_));
 sg13g2_o21ai_1 _6153_ (.B1(net453),
    .Y(_2777_),
    .A1(_2771_),
    .A2(_2775_));
 sg13g2_a21oi_1 _6154_ (.A1(_2771_),
    .A2(_2775_),
    .Y(_0433_),
    .B1(_2777_));
 sg13g2_a21o_1 _6155_ (.A2(_2776_),
    .A1(_2770_),
    .B1(_2774_),
    .X(_2778_));
 sg13g2_o21ai_1 _6156_ (.B1(_2772_),
    .Y(_2779_),
    .A1(net511),
    .A2(_0621_));
 sg13g2_nor2_1 _6157_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][8] ),
    .B(_2779_),
    .Y(_2780_));
 sg13g2_xor2_1 _6158_ (.B(_2779_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][8] ),
    .X(_2781_));
 sg13g2_nand2b_1 _6159_ (.Y(_2782_),
    .B(net1425),
    .A_N(_2781_));
 sg13g2_inv_1 _6160_ (.Y(_2783_),
    .A(_2782_));
 sg13g2_xnor2_1 _6161_ (.Y(_2784_),
    .A(net1425),
    .B(_2781_));
 sg13g2_o21ai_1 _6162_ (.B1(net453),
    .Y(_2785_),
    .A1(_2778_),
    .A2(_2784_));
 sg13g2_a21oi_1 _6163_ (.A1(_2778_),
    .A2(net1426),
    .Y(_0434_),
    .B1(_2785_));
 sg13g2_a21o_1 _6164_ (.A2(_2784_),
    .A1(_2778_),
    .B1(_2783_),
    .X(_2786_));
 sg13g2_nor2_1 _6165_ (.A(net507),
    .B(_2780_),
    .Y(_2787_));
 sg13g2_xnor2_1 _6166_ (.Y(_2788_),
    .A(net1371),
    .B(_2787_));
 sg13g2_and2_1 _6167_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[7] ),
    .B(_2788_),
    .X(_2789_));
 sg13g2_xnor2_1 _6168_ (.Y(_2790_),
    .A(_0622_),
    .B(_2788_));
 sg13g2_nor2_1 _6169_ (.A(_2786_),
    .B(_2790_),
    .Y(_2791_));
 sg13g2_a21oi_1 _6170_ (.A1(_2786_),
    .A2(_2790_),
    .Y(_2792_),
    .B1(net424));
 sg13g2_nor2b_1 _6171_ (.A(_2791_),
    .B_N(_2792_),
    .Y(_0435_));
 sg13g2_a21o_1 _6172_ (.A2(_2790_),
    .A1(_2786_),
    .B1(_2789_),
    .X(_2793_));
 sg13g2_a21oi_1 _6173_ (.A1(_0623_),
    .A2(_2780_),
    .Y(_2794_),
    .B1(net507));
 sg13g2_nor2_1 _6174_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][10] ),
    .B(_2794_),
    .Y(_2795_));
 sg13g2_xnor2_1 _6175_ (.Y(_2796_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][10] ),
    .B(_2794_));
 sg13g2_and2_1 _6176_ (.A(net1491),
    .B(_2796_),
    .X(_2797_));
 sg13g2_xor2_1 _6177_ (.B(_2796_),
    .A(net1491),
    .X(_2798_));
 sg13g2_o21ai_1 _6178_ (.B1(net454),
    .Y(_2799_),
    .A1(_2793_),
    .A2(_2798_));
 sg13g2_a21oi_1 _6179_ (.A1(_2793_),
    .A2(_2798_),
    .Y(_0436_),
    .B1(_2799_));
 sg13g2_a21o_2 _6180_ (.A2(_2798_),
    .A1(_2793_),
    .B1(_2797_),
    .X(_2800_));
 sg13g2_nor2_1 _6181_ (.A(net510),
    .B(_2795_),
    .Y(_2801_));
 sg13g2_xnor2_1 _6182_ (.Y(_2802_),
    .A(net1130),
    .B(_2801_));
 sg13g2_and2_1 _6183_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[9] ),
    .B(_2802_),
    .X(_2803_));
 sg13g2_xor2_1 _6184_ (.B(_2802_),
    .A(net1508),
    .X(_2804_));
 sg13g2_nor2_1 _6185_ (.A(_2800_),
    .B(_2804_),
    .Y(_2805_));
 sg13g2_a21oi_1 _6186_ (.A1(_2800_),
    .A2(_2804_),
    .Y(_2806_),
    .B1(net424));
 sg13g2_nor2b_1 _6187_ (.A(_2805_),
    .B_N(_2806_),
    .Y(_0437_));
 sg13g2_a21oi_1 _6188_ (.A1(_2800_),
    .A2(_2804_),
    .Y(_2807_),
    .B1(_2803_));
 sg13g2_a21o_1 _6189_ (.A2(_2804_),
    .A1(_2800_),
    .B1(_2803_),
    .X(_2808_));
 sg13g2_a21oi_1 _6190_ (.A1(_0624_),
    .A2(_2795_),
    .Y(_2809_),
    .B1(net510));
 sg13g2_xnor2_1 _6191_ (.Y(_2810_),
    .A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][12] ),
    .B(_2809_));
 sg13g2_and2_1 _6192_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[10] ),
    .B(_2810_),
    .X(_2811_));
 sg13g2_xnor2_1 _6193_ (.Y(_2812_),
    .A(net1343),
    .B(_2810_));
 sg13g2_inv_1 _6194_ (.Y(_2813_),
    .A(_2812_));
 sg13g2_o21ai_1 _6195_ (.B1(net454),
    .Y(_2814_),
    .A1(_2807_),
    .A2(_2812_));
 sg13g2_a21oi_1 _6196_ (.A1(_2807_),
    .A2(net1344),
    .Y(_0438_),
    .B1(_2814_));
 sg13g2_a21oi_1 _6197_ (.A1(_2808_),
    .A2(_2813_),
    .Y(_2815_),
    .B1(_2811_));
 sg13g2_mux2_1 _6198_ (.A0(_2809_),
    .A1(net510),
    .S(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][12] ),
    .X(_2816_));
 sg13g2_xor2_1 _6199_ (.B(_2816_),
    .A(net1281),
    .X(_2817_));
 sg13g2_o21ai_1 _6200_ (.B1(net454),
    .Y(_2818_),
    .A1(_2815_),
    .A2(_2817_));
 sg13g2_a21oi_1 _6201_ (.A1(_2815_),
    .A2(net1282),
    .Y(_0439_),
    .B1(_2818_));
 sg13g2_and2_1 _6202_ (.A(net466),
    .B(net761),
    .X(_0440_));
 sg13g2_nor2_1 _6203_ (.A(net759),
    .B(net426),
    .Y(_0441_));
 sg13g2_nand2_1 _6204_ (.Y(_2819_),
    .A(net1005),
    .B(net508));
 sg13g2_xor2_1 _6205_ (.B(net508),
    .A(net1005),
    .X(_2820_));
 sg13g2_nand2_1 _6206_ (.Y(_2821_),
    .A(net759),
    .B(_2820_));
 sg13g2_o21ai_1 _6207_ (.B1(net466),
    .Y(_2822_),
    .A1(net759),
    .A2(_2820_));
 sg13g2_nor2b_1 _6208_ (.A(_2822_),
    .B_N(_2821_),
    .Y(_0442_));
 sg13g2_xnor2_1 _6209_ (.Y(_2823_),
    .A(net508),
    .B(net1049));
 sg13g2_and3_1 _6210_ (.X(_2824_),
    .A(_2819_),
    .B(_2821_),
    .C(_2823_));
 sg13g2_a21oi_1 _6211_ (.A1(_2819_),
    .A2(_2821_),
    .Y(_2825_),
    .B1(_2823_));
 sg13g2_nor3_1 _6212_ (.A(net426),
    .B(_2824_),
    .C(_2825_),
    .Y(_0443_));
 sg13g2_a21oi_1 _6213_ (.A1(net508),
    .A2(net1049),
    .Y(_2826_),
    .B1(_2825_));
 sg13g2_nand2_1 _6214_ (.Y(_2827_),
    .A(net417),
    .B(net1329));
 sg13g2_xor2_1 _6215_ (.B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][4] ),
    .A(net508),
    .X(_2828_));
 sg13g2_or2_1 _6216_ (.X(_2829_),
    .B(_2828_),
    .A(_2826_));
 sg13g2_nand2_1 _6217_ (.Y(_2830_),
    .A(net462),
    .B(_2829_));
 sg13g2_a21oi_1 _6218_ (.A1(_2826_),
    .A2(_2828_),
    .Y(_0444_),
    .B1(_2830_));
 sg13g2_nand2_1 _6219_ (.Y(_2831_),
    .A(net508),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][5] ));
 sg13g2_xnor2_1 _6220_ (.Y(_2832_),
    .A(net509),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][5] ));
 sg13g2_nand3_1 _6221_ (.B(_2829_),
    .C(_2832_),
    .A(_2827_),
    .Y(_2833_));
 sg13g2_a21o_1 _6222_ (.A2(_2829_),
    .A1(_2827_),
    .B1(_2832_),
    .X(_2834_));
 sg13g2_and3_1 _6223_ (.X(_0445_),
    .A(net455),
    .B(net1330),
    .C(_2834_));
 sg13g2_and2_1 _6224_ (.A(_2831_),
    .B(_2834_),
    .X(_2835_));
 sg13g2_nor2_1 _6225_ (.A(net417),
    .B(net1235),
    .Y(_2836_));
 sg13g2_nand2_1 _6226_ (.Y(_2837_),
    .A(net417),
    .B(net1235));
 sg13g2_nand2b_1 _6227_ (.Y(_2838_),
    .B(_2837_),
    .A_N(_2836_));
 sg13g2_o21ai_1 _6228_ (.B1(net454),
    .Y(_2839_),
    .A1(_2835_),
    .A2(_2838_));
 sg13g2_a21oi_1 _6229_ (.A1(_2835_),
    .A2(_2838_),
    .Y(_0446_),
    .B1(_2839_));
 sg13g2_xnor2_1 _6230_ (.Y(_2840_),
    .A(net509),
    .B(net1267));
 sg13g2_o21ai_1 _6231_ (.B1(_2837_),
    .Y(_2841_),
    .A1(_2835_),
    .A2(_2836_));
 sg13g2_and2_1 _6232_ (.A(_2840_),
    .B(_2841_),
    .X(_2842_));
 sg13g2_o21ai_1 _6233_ (.B1(net455),
    .Y(_2843_),
    .A1(_2840_),
    .A2(_2841_));
 sg13g2_nor2_1 _6234_ (.A(_2842_),
    .B(_2843_),
    .Y(_0447_));
 sg13g2_a21oi_1 _6235_ (.A1(net417),
    .A2(net1267),
    .Y(_2844_),
    .B1(_2842_));
 sg13g2_xnor2_1 _6236_ (.Y(_2845_),
    .A(net508),
    .B(net1071));
 sg13g2_nor2_1 _6237_ (.A(_2844_),
    .B(_2845_),
    .Y(_2846_));
 sg13g2_a21oi_1 _6238_ (.A1(_2844_),
    .A2(_2845_),
    .Y(_2847_),
    .B1(net424));
 sg13g2_nor2b_1 _6239_ (.A(_2846_),
    .B_N(_2847_),
    .Y(_0448_));
 sg13g2_a21oi_1 _6240_ (.A1(net508),
    .A2(net1071),
    .Y(_2848_),
    .B1(_2846_));
 sg13g2_xor2_1 _6241_ (.B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][9] ),
    .A(net510),
    .X(_2849_));
 sg13g2_or2_1 _6242_ (.X(_2850_),
    .B(_2849_),
    .A(_2848_));
 sg13g2_nand2_1 _6243_ (.Y(_2851_),
    .A(net455),
    .B(_2850_));
 sg13g2_a21oi_1 _6244_ (.A1(net1072),
    .A2(_2849_),
    .Y(_0449_),
    .B1(_2851_));
 sg13g2_o21ai_1 _6245_ (.B1(_2850_),
    .Y(_2852_),
    .A1(net510),
    .A2(_0563_));
 sg13g2_xnor2_1 _6246_ (.Y(_2853_),
    .A(net510),
    .B(net1099));
 sg13g2_o21ai_1 _6247_ (.B1(net455),
    .Y(_2854_),
    .A1(_2852_),
    .A2(_2853_));
 sg13g2_a21oi_1 _6248_ (.A1(_2852_),
    .A2(_2853_),
    .Y(_0450_),
    .B1(_2854_));
 sg13g2_nand2b_1 _6249_ (.Y(_2855_),
    .B(_2853_),
    .A_N(_2850_));
 sg13g2_o21ai_1 _6250_ (.B1(net417),
    .Y(_2856_),
    .A1(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][9] ),
    .A2(net1099));
 sg13g2_and3_1 _6251_ (.X(_0451_),
    .A(net455),
    .B(_2855_),
    .C(net1100));
 sg13g2_nand2b_1 _6252_ (.Y(_2857_),
    .B(net1041),
    .A_N(net967));
 sg13g2_nand2_1 _6253_ (.Y(_2858_),
    .A(net967),
    .B(_0543_));
 sg13g2_a21oi_1 _6254_ (.A1(net402),
    .A2(net968),
    .Y(_0452_),
    .B1(net421));
 sg13g2_nand2_1 _6255_ (.Y(_2859_),
    .A(net967),
    .B(_0605_));
 sg13g2_a21o_2 _6256_ (.A2(_2859_),
    .A1(net402),
    .B1(net555),
    .X(_2860_));
 sg13g2_nand3_1 _6257_ (.B(net402),
    .C(_2859_),
    .A(net555),
    .Y(_2861_));
 sg13g2_a21oi_1 _6258_ (.A1(_2860_),
    .A2(_2861_),
    .Y(_0453_),
    .B1(net421));
 sg13g2_nand2_2 _6259_ (.Y(_2862_),
    .A(net506),
    .B(net555));
 sg13g2_a21oi_1 _6260_ (.A1(_2860_),
    .A2(_2862_),
    .Y(_0454_),
    .B1(net421));
 sg13g2_nor2_1 _6261_ (.A(net967),
    .B(net555),
    .Y(_2863_));
 sg13g2_nor3_1 _6262_ (.A(net506),
    .B(net1070),
    .C(_2863_),
    .Y(_2864_));
 sg13g2_o21ai_1 _6263_ (.B1(net1070),
    .Y(_2865_),
    .A1(net506),
    .A2(_2863_));
 sg13g2_nor2b_1 _6264_ (.A(_2864_),
    .B_N(_2865_),
    .Y(_2866_));
 sg13g2_o21ai_1 _6265_ (.B1(net1041),
    .Y(_2867_),
    .A1(net967),
    .A2(net555));
 sg13g2_and2_1 _6266_ (.A(net444),
    .B(_2867_),
    .X(_2868_));
 sg13g2_nor2_1 _6267_ (.A(net421),
    .B(_2867_),
    .Y(_2869_));
 sg13g2_mux2_1 _6268_ (.A0(_2868_),
    .A1(_2869_),
    .S(_2866_),
    .X(_0458_));
 sg13g2_o21ai_1 _6269_ (.B1(net1070),
    .Y(_2870_),
    .A1(_0543_),
    .A2(net939));
 sg13g2_nand3b_1 _6270_ (.B(net1041),
    .C(_0605_),
    .Y(_2871_),
    .A_N(net1070));
 sg13g2_and2_1 _6271_ (.A(_2870_),
    .B(_2871_),
    .X(_2872_));
 sg13g2_nor2_2 _6272_ (.A(_2867_),
    .B(_2872_),
    .Y(_2873_));
 sg13g2_nor2_1 _6273_ (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[0].y_shr[0] ),
    .B(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[0].y_shr[11] ),
    .Y(_2874_));
 sg13g2_nor3_1 _6274_ (.A(net506),
    .B(net555),
    .C(_2874_),
    .Y(_2875_));
 sg13g2_a21o_1 _6275_ (.A2(net555),
    .A1(net506),
    .B1(_2875_),
    .X(_2876_));
 sg13g2_xnor2_1 _6276_ (.Y(_2877_),
    .A(_0543_),
    .B(_2876_));
 sg13g2_o21ai_1 _6277_ (.B1(net444),
    .Y(_2878_),
    .A1(_2873_),
    .A2(_2877_));
 sg13g2_a21oi_1 _6278_ (.A1(_2873_),
    .A2(_2877_),
    .Y(_0459_),
    .B1(_2878_));
 sg13g2_a21oi_1 _6279_ (.A1(net939),
    .A2(net1070),
    .Y(_2879_),
    .B1(_2864_));
 sg13g2_a221oi_1 _6280_ (.B2(net1041),
    .C1(_2864_),
    .B1(_2876_),
    .A1(net939),
    .Y(_2880_),
    .A2(net1070));
 sg13g2_nor3_1 _6281_ (.A(net421),
    .B(_2873_),
    .C(_2880_),
    .Y(_0460_));
 sg13g2_nor2b_1 _6282_ (.A(_2879_),
    .B_N(_2868_),
    .Y(_0461_));
 sg13g2_nand2_2 _6283_ (.Y(_2881_),
    .A(net1041),
    .B(net506));
 sg13g2_nand2_2 _6284_ (.Y(_2882_),
    .A(net1043),
    .B(_2881_));
 sg13g2_xnor2_1 _6285_ (.Y(_2883_),
    .A(net1043),
    .B(_2881_));
 sg13g2_nand2b_1 _6286_ (.Y(_2884_),
    .B(_2883_),
    .A_N(net402));
 sg13g2_nand2b_1 _6287_ (.Y(_2885_),
    .B(net402),
    .A_N(_2883_));
 sg13g2_and3_1 _6288_ (.X(_0465_),
    .A(net444),
    .B(_2884_),
    .C(_2885_));
 sg13g2_o21ai_1 _6289_ (.B1(net444),
    .Y(_2886_),
    .A1(net555),
    .A2(_2881_));
 sg13g2_a21oi_1 _6290_ (.A1(net402),
    .A2(_2882_),
    .Y(_0466_),
    .B1(_2886_));
 sg13g2_nand2_1 _6291_ (.Y(_2887_),
    .A(_2882_),
    .B(_2885_));
 sg13g2_nor2_1 _6292_ (.A(_2872_),
    .B(_2887_),
    .Y(_2888_));
 sg13g2_nand2_1 _6293_ (.Y(_2889_),
    .A(_2872_),
    .B(_2887_));
 sg13g2_nand2_1 _6294_ (.Y(_2890_),
    .A(net444),
    .B(_2889_));
 sg13g2_nor2_1 _6295_ (.A(_2888_),
    .B(_2890_),
    .Y(_0470_));
 sg13g2_nand3_1 _6296_ (.B(_2883_),
    .C(_2889_),
    .A(_2870_),
    .Y(_2891_));
 sg13g2_a21o_1 _6297_ (.A2(_2889_),
    .A1(_2870_),
    .B1(_2883_),
    .X(_2892_));
 sg13g2_and3_1 _6298_ (.X(_0471_),
    .A(net444),
    .B(_2891_),
    .C(_2892_));
 sg13g2_nor2b_1 _6299_ (.A(_2872_),
    .B_N(_2882_),
    .Y(_2893_));
 sg13g2_a21oi_1 _6300_ (.A1(_2892_),
    .A2(_2893_),
    .Y(_0472_),
    .B1(_2890_));
 sg13g2_nand2_1 _6301_ (.Y(_2894_),
    .A(net444),
    .B(_2871_));
 sg13g2_a21oi_1 _6302_ (.A1(_2870_),
    .A2(_2887_),
    .Y(_0473_),
    .B1(_2894_));
 sg13g2_and2_1 _6303_ (.A(net462),
    .B(net765),
    .X(_0477_));
 sg13g2_and2_1 _6304_ (.A(net462),
    .B(net767),
    .X(_0478_));
 sg13g2_and2_1 _6305_ (.A(net462),
    .B(net764),
    .X(_0479_));
 sg13g2_and2_1 _6306_ (.A(net462),
    .B(net769),
    .X(_0480_));
 sg13g2_and2_1 _6307_ (.A(net454),
    .B(net786),
    .X(_0481_));
 sg13g2_and2_1 _6308_ (.A(net446),
    .B(net775),
    .X(_0482_));
 sg13g2_and2_1 _6309_ (.A(net446),
    .B(net787),
    .X(_0483_));
 sg13g2_and2_1 _6310_ (.A(net446),
    .B(net778),
    .X(_0484_));
 sg13g2_and2_1 _6311_ (.A(net446),
    .B(net780),
    .X(_0485_));
 sg13g2_nor2_1 _6312_ (.A(net758),
    .B(net422),
    .Y(_0486_));
 sg13g2_xnor2_1 _6313_ (.Y(_2895_),
    .A(net506),
    .B(net815));
 sg13g2_nor2_1 _6314_ (.A(net758),
    .B(_2895_),
    .Y(_2896_));
 sg13g2_a21o_1 _6315_ (.A2(_2895_),
    .A1(net758),
    .B1(net422),
    .X(_2897_));
 sg13g2_nor2_1 _6316_ (.A(_2896_),
    .B(_2897_),
    .Y(_0487_));
 sg13g2_a21oi_1 _6317_ (.A1(_0605_),
    .A2(net815),
    .Y(_0488_),
    .B1(_2897_));
 sg13g2_and2_1 _6318_ (.A(net465),
    .B(net806),
    .X(_0489_));
 sg13g2_and2_1 _6319_ (.A(net465),
    .B(net802),
    .X(_0490_));
 sg13g2_and2_1 _6320_ (.A(net464),
    .B(net779),
    .X(_0491_));
 sg13g2_and2_1 _6321_ (.A(net463),
    .B(net784),
    .X(_0492_));
 sg13g2_and2_1 _6322_ (.A(net464),
    .B(net793),
    .X(_0493_));
 sg13g2_and2_1 _6323_ (.A(net468),
    .B(net801),
    .X(_0494_));
 sg13g2_and2_1 _6324_ (.A(net462),
    .B(net771),
    .X(_0495_));
 sg13g2_and2_1 _6325_ (.A(net466),
    .B(net796),
    .X(_0496_));
 sg13g2_and2_1 _6326_ (.A(net462),
    .B(net785),
    .X(_0497_));
 sg13g2_and2_1 _6327_ (.A(net462),
    .B(net794),
    .X(_0498_));
 sg13g2_and2_1 _6328_ (.A(net463),
    .B(net789),
    .X(_0499_));
 sg13g2_and2_1 _6329_ (.A(net469),
    .B(net839),
    .X(_0500_));
 sg13g2_nor2_1 _6330_ (.A(net763),
    .B(net374),
    .Y(_0501_));
 sg13g2_and2_1 _6331_ (.A(net763),
    .B(net1007),
    .X(_2898_));
 sg13g2_nor3_1 _6332_ (.A(_0958_),
    .B(net374),
    .C(_2898_),
    .Y(_0502_));
 sg13g2_and2_1 _6333_ (.A(net898),
    .B(_2898_),
    .X(_2899_));
 sg13g2_nor2_1 _6334_ (.A(net898),
    .B(_2898_),
    .Y(_2900_));
 sg13g2_nor3_1 _6335_ (.A(net374),
    .B(_2899_),
    .C(net899),
    .Y(_0503_));
 sg13g2_and2_1 _6336_ (.A(net931),
    .B(_2899_),
    .X(_2901_));
 sg13g2_nor2_1 _6337_ (.A(net931),
    .B(_2899_),
    .Y(_2902_));
 sg13g2_nor3_1 _6338_ (.A(net374),
    .B(_2901_),
    .C(net932),
    .Y(_0504_));
 sg13g2_and2_1 _6339_ (.A(net926),
    .B(_2901_),
    .X(_2903_));
 sg13g2_nor2_1 _6340_ (.A(net926),
    .B(_2901_),
    .Y(_2904_));
 sg13g2_nor3_1 _6341_ (.A(net374),
    .B(_2903_),
    .C(net927),
    .Y(_0505_));
 sg13g2_o21ai_1 _6342_ (.B1(net378),
    .Y(_2905_),
    .A1(net844),
    .A2(_2903_));
 sg13g2_a21oi_1 _6343_ (.A1(net844),
    .A2(_2903_),
    .Y(_0506_),
    .B1(_2905_));
 sg13g2_nand3_1 _6344_ (.B(net1114),
    .C(_2903_),
    .A(net844),
    .Y(_2906_));
 sg13g2_a21o_1 _6345_ (.A2(_2903_),
    .A1(net844),
    .B1(net1114),
    .X(_2907_));
 sg13g2_and3_1 _6346_ (.X(_0507_),
    .A(net378),
    .B(_2906_),
    .C(_2907_));
 sg13g2_nor2_1 _6347_ (.A(_0547_),
    .B(_2906_),
    .Y(_2908_));
 sg13g2_and2_1 _6348_ (.A(_0547_),
    .B(_2906_),
    .X(_2909_));
 sg13g2_nor3_1 _6349_ (.A(net374),
    .B(_2908_),
    .C(net1108),
    .Y(_0508_));
 sg13g2_and2_1 _6350_ (.A(net956),
    .B(_2908_),
    .X(_2910_));
 sg13g2_nor2_1 _6351_ (.A(net956),
    .B(_2908_),
    .Y(_2911_));
 sg13g2_nor3_1 _6352_ (.A(net374),
    .B(_2910_),
    .C(net957),
    .Y(_0509_));
 sg13g2_o21ai_1 _6353_ (.B1(net378),
    .Y(_2912_),
    .A1(net847),
    .A2(_2910_));
 sg13g2_a21oi_1 _6354_ (.A1(net847),
    .A2(_2910_),
    .Y(_0510_),
    .B1(_2912_));
 sg13g2_and3_1 _6355_ (.X(_2913_),
    .A(net847),
    .B(net880),
    .C(_2910_));
 sg13g2_a21oi_1 _6356_ (.A1(net847),
    .A2(_2910_),
    .Y(_2914_),
    .B1(net880));
 sg13g2_nor3_1 _6357_ (.A(net374),
    .B(_2913_),
    .C(net881),
    .Y(_0511_));
 sg13g2_and2_1 _6358_ (.A(net975),
    .B(_2913_),
    .X(_2915_));
 sg13g2_nor2_1 _6359_ (.A(net975),
    .B(_2913_),
    .Y(_2916_));
 sg13g2_nor3_1 _6360_ (.A(net375),
    .B(_2915_),
    .C(_2916_),
    .Y(_0512_));
 sg13g2_and2_1 _6361_ (.A(net981),
    .B(_2915_),
    .X(_2917_));
 sg13g2_nor2_1 _6362_ (.A(net981),
    .B(_2915_),
    .Y(_2918_));
 sg13g2_nor3_1 _6363_ (.A(net375),
    .B(_2917_),
    .C(_2918_),
    .Y(_0513_));
 sg13g2_and2_1 _6364_ (.A(net958),
    .B(_2917_),
    .X(_2919_));
 sg13g2_nor2_1 _6365_ (.A(net958),
    .B(_2917_),
    .Y(_2920_));
 sg13g2_nor3_1 _6366_ (.A(net375),
    .B(_2919_),
    .C(net959),
    .Y(_0514_));
 sg13g2_and2_1 _6367_ (.A(net1022),
    .B(_2919_),
    .X(_2921_));
 sg13g2_o21ai_1 _6368_ (.B1(net377),
    .Y(_2922_),
    .A1(net1022),
    .A2(_2919_));
 sg13g2_nor2_1 _6369_ (.A(_2921_),
    .B(_2922_),
    .Y(_0515_));
 sg13g2_o21ai_1 _6370_ (.B1(net377),
    .Y(_2923_),
    .A1(net854),
    .A2(_2921_));
 sg13g2_a21oi_1 _6371_ (.A1(net854),
    .A2(_2921_),
    .Y(_0516_),
    .B1(_2923_));
 sg13g2_a21oi_1 _6372_ (.A1(net854),
    .A2(_2921_),
    .Y(_2924_),
    .B1(net916));
 sg13g2_and3_1 _6373_ (.X(_2925_),
    .A(net854),
    .B(net916),
    .C(_2921_));
 sg13g2_nor3_1 _6374_ (.A(net375),
    .B(net917),
    .C(_2925_),
    .Y(_0517_));
 sg13g2_a21oi_1 _6375_ (.A1(net1029),
    .A2(_2925_),
    .Y(_2926_),
    .B1(net375));
 sg13g2_o21ai_1 _6376_ (.B1(_2926_),
    .Y(_2927_),
    .A1(net1029),
    .A2(_2925_));
 sg13g2_inv_1 _6377_ (.Y(_0518_),
    .A(_2927_));
 sg13g2_and2_1 _6378_ (.A(net878),
    .B(net442),
    .X(_0521_));
 sg13g2_a21oi_1 _6379_ (.A1(_2860_),
    .A2(_2862_),
    .Y(_0455_),
    .B1(net421));
 sg13g2_a21oi_1 _6380_ (.A1(_2860_),
    .A2(_2862_),
    .Y(_0456_),
    .B1(net421));
 sg13g2_a21oi_1 _6381_ (.A1(_2860_),
    .A2(_2862_),
    .Y(_0457_),
    .B1(net421));
 sg13g2_a21oi_1 _6382_ (.A1(_2873_),
    .A2(_2877_),
    .Y(_0462_),
    .B1(_2878_));
 sg13g2_nor3_1 _6383_ (.A(net422),
    .B(_2873_),
    .C(_2880_),
    .Y(_0463_));
 sg13g2_nor2b_1 _6384_ (.A(_2879_),
    .B_N(_2868_),
    .Y(_0464_));
 sg13g2_a21oi_1 _6385_ (.A1(net402),
    .A2(_2882_),
    .Y(_0467_),
    .B1(_2886_));
 sg13g2_a21oi_1 _6386_ (.A1(net402),
    .A2(_2882_),
    .Y(_0468_),
    .B1(_2886_));
 sg13g2_a21oi_1 _6387_ (.A1(_2857_),
    .A2(_2882_),
    .Y(_0469_),
    .B1(_2886_));
 sg13g2_and3_1 _6388_ (.X(_0474_),
    .A(net447),
    .B(_2891_),
    .C(_2892_));
 sg13g2_a21oi_1 _6389_ (.A1(_2892_),
    .A2(_2893_),
    .Y(_0475_),
    .B1(_2890_));
 sg13g2_a21oi_1 _6390_ (.A1(_2870_),
    .A2(_2887_),
    .Y(_0476_),
    .B1(_2894_));
 sg13g2_dfrbpq_2 _6391_ (.RESET_B(net725),
    .D(_0000_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[0].y_shr[11] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _6392_ (.RESET_B(net574),
    .D(_0001_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[0].y_shr[10] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _6393_ (.RESET_B(net573),
    .D(net861),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[0].y_shr[0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _6394_ (.RESET_B(net572),
    .D(net823),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[0][0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6395_ (.RESET_B(net571),
    .D(net930),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[5] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6396_ (.RESET_B(net569),
    .D(net836),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[9] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6397_ (.RESET_B(net567),
    .D(net814),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[10] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6398_ (.RESET_B(net565),
    .D(_0007_),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.clk_div_cnt[0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6399_ (.RESET_B(net564),
    .D(_0008_),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.clk_div_cnt[1] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _6400_ (.RESET_B(net563),
    .D(net897),
    .Q(net21),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6401_ (.RESET_B(net561),
    .D(net1067),
    .Q(net22),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6402_ (.RESET_B(net559),
    .D(_0011_),
    .Q(pwm_data),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6403_ (.RESET_B(net558),
    .D(net884),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6404_ (.RESET_B(net556),
    .D(net908),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[1] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6405_ (.RESET_B(net370),
    .D(net894),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[2] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6406_ (.RESET_B(net368),
    .D(net911),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6407_ (.RESET_B(net366),
    .D(net945),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[4] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6408_ (.RESET_B(net364),
    .D(net868),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[6] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6409_ (.RESET_B(net362),
    .D(net871),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _6410_ (.RESET_B(net360),
    .D(net891),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[8] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6411_ (.RESET_B(net358),
    .D(net858),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[0] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6412_ (.RESET_B(net356),
    .D(net876),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[1] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6413_ (.RESET_B(net354),
    .D(_0022_),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[2] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_1 _6414_ (.RESET_B(net352),
    .D(net938),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[3] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _6415_ (.RESET_B(net350),
    .D(_0024_),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[4] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _6416_ (.RESET_B(net348),
    .D(_0025_),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[5] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _6417_ (.RESET_B(net346),
    .D(net1032),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[6] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _6418_ (.RESET_B(net344),
    .D(net1021),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _6419_ (.RESET_B(net342),
    .D(net843),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[8] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6420_ (.RESET_B(net340),
    .D(_0029_),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[9] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6421_ (.RESET_B(net338),
    .D(net984),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[10] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _6422_ (.RESET_B(net336),
    .D(_0031_),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _6423_ (.RESET_B(net334),
    .D(net1025),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _6424_ (.RESET_B(net332),
    .D(net921),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _6425_ (.RESET_B(net330),
    .D(net979),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[3] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _6426_ (.RESET_B(net328),
    .D(_0035_),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[4] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _6427_ (.RESET_B(net326),
    .D(_0036_),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _6428_ (.RESET_B(net324),
    .D(net943),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[6] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _6429_ (.RESET_B(net322),
    .D(net902),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _6430_ (.RESET_B(net320),
    .D(_0039_),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[8] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _6431_ (.RESET_B(net318),
    .D(net1002),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[9] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _6432_ (.RESET_B(net316),
    .D(net864),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[10] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _6433_ (.RESET_B(net314),
    .D(_0042_),
    .Q(\u_angle_cordic_12b_pmod.u_vga_top.pixel_clk_en ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_1 _6434_ (.RESET_B(net313),
    .D(_0043_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[0] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6435_ (.RESET_B(net312),
    .D(_0044_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6436_ (.RESET_B(net311),
    .D(_0045_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6437_ (.RESET_B(net310),
    .D(_0046_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6438_ (.RESET_B(net309),
    .D(_0047_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[4] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6439_ (.RESET_B(net308),
    .D(_0048_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[5] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6440_ (.RESET_B(net307),
    .D(net782),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[6] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6441_ (.RESET_B(net306),
    .D(net777),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[7] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6442_ (.RESET_B(net305),
    .D(_0051_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[8] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6443_ (.RESET_B(net304),
    .D(_0052_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[9] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6444_ (.RESET_B(net303),
    .D(_0053_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[10] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6445_ (.RESET_B(net302),
    .D(_0054_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.COSout[11] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6446_ (.RESET_B(net301),
    .D(net1180),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.up ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6447_ (.RESET_B(net299),
    .D(_0056_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6448_ (.RESET_B(net297),
    .D(net925),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6449_ (.RESET_B(net295),
    .D(_0058_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[2] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6450_ (.RESET_B(net293),
    .D(net955),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[3] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6451_ (.RESET_B(net291),
    .D(net949),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[4] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _6452_ (.RESET_B(net289),
    .D(_0061_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[5] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6453_ (.RESET_B(net287),
    .D(net953),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[6] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6454_ (.RESET_B(net285),
    .D(net886),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[7] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6455_ (.RESET_B(net283),
    .D(_0064_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _6456_ (.RESET_B(net281),
    .D(net1013),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[9] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _6457_ (.RESET_B(net279),
    .D(_0066_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[10] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6458_ (.RESET_B(net277),
    .D(_0067_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[11] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _6459_ (.RESET_B(net275),
    .D(_0068_),
    .Q(\u_angle_cordic_12b_pmod.waveform_sel_reg[0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6460_ (.RESET_B(net274),
    .D(_0069_),
    .Q(\u_angle_cordic_12b_pmod.waveform_sel_reg[1] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _6461_ (.RESET_B(net273),
    .D(_0070_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _6462_ (.RESET_B(net271),
    .D(_0071_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[1] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6463_ (.RESET_B(net269),
    .D(_0072_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[2] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _6464_ (.RESET_B(net267),
    .D(_0073_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6465_ (.RESET_B(net265),
    .D(_0074_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[4] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6466_ (.RESET_B(net263),
    .D(_0075_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[5] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6467_ (.RESET_B(net261),
    .D(_0076_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[6] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6468_ (.RESET_B(net259),
    .D(net829),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6469_ (.RESET_B(net257),
    .D(_0078_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[8] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _6470_ (.RESET_B(net255),
    .D(_0079_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[9] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _6471_ (.RESET_B(net253),
    .D(_0080_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[10] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _6472_ (.RESET_B(net251),
    .D(_0081_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[11] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6473_ (.RESET_B(net249),
    .D(_0082_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp[11] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _6474_ (.RESET_B(net248),
    .D(_0083_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6475_ (.RESET_B(net247),
    .D(_0084_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6476_ (.RESET_B(net246),
    .D(_0085_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][2] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6477_ (.RESET_B(net245),
    .D(net1059),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][3] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6478_ (.RESET_B(net244),
    .D(_0087_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][4] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6479_ (.RESET_B(net243),
    .D(net1061),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][5] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6480_ (.RESET_B(net242),
    .D(_0089_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][6] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6481_ (.RESET_B(net241),
    .D(net1176),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][7] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6482_ (.RESET_B(net240),
    .D(net1152),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][8] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6483_ (.RESET_B(net239),
    .D(net1116),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][9] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6484_ (.RESET_B(net238),
    .D(_0093_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][10] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _6485_ (.RESET_B(net237),
    .D(_0094_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].z_sign ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6486_ (.RESET_B(net236),
    .D(_0095_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6487_ (.RESET_B(net235),
    .D(net1105),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][1] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6488_ (.RESET_B(net234),
    .D(net1357),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][2] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _6489_ (.RESET_B(net233),
    .D(_0098_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][3] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _6490_ (.RESET_B(net232),
    .D(_0099_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][4] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _6491_ (.RESET_B(net231),
    .D(_0100_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][5] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6492_ (.RESET_B(net230),
    .D(_0101_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][6] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _6493_ (.RESET_B(net229),
    .D(_0102_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _6494_ (.RESET_B(net228),
    .D(_0103_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[1] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _6495_ (.RESET_B(net227),
    .D(net1184),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[2] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _6496_ (.RESET_B(net226),
    .D(_0105_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[3] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _6497_ (.RESET_B(net225),
    .D(net1301),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[4] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6498_ (.RESET_B(net224),
    .D(net1310),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[10] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6499_ (.RESET_B(net223),
    .D(net964),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6500_ (.RESET_B(net222),
    .D(net992),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][1] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6501_ (.RESET_B(net221),
    .D(_0110_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][2] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6502_ (.RESET_B(net220),
    .D(_0111_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][3] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6503_ (.RESET_B(net219),
    .D(_0112_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][4] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6504_ (.RESET_B(net218),
    .D(net1405),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][5] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6505_ (.RESET_B(net217),
    .D(_0114_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][6] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _6506_ (.RESET_B(net216),
    .D(_0115_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][7] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _6507_ (.RESET_B(net215),
    .D(_0116_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][8] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _6508_ (.RESET_B(net214),
    .D(net1513),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][9] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _6509_ (.RESET_B(net213),
    .D(net1529),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][10] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _6510_ (.RESET_B(net212),
    .D(net1362),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][11] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _6511_ (.RESET_B(net211),
    .D(net1200),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][12] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6512_ (.RESET_B(net210),
    .D(_0121_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6513_ (.RESET_B(net209),
    .D(_0122_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6514_ (.RESET_B(net208),
    .D(net1028),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][2] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6515_ (.RESET_B(net207),
    .D(_0124_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][3] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6516_ (.RESET_B(net206),
    .D(net1081),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][4] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6517_ (.RESET_B(net205),
    .D(_0126_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][5] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6518_ (.RESET_B(net204),
    .D(net1193),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][6] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6519_ (.RESET_B(net203),
    .D(net1141),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][7] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6520_ (.RESET_B(net202),
    .D(net1111),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][8] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6521_ (.RESET_B(net201),
    .D(_0130_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][9] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6522_ (.RESET_B(net200),
    .D(_0131_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][10] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _6523_ (.RESET_B(net199),
    .D(net819),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].z_sign ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _6524_ (.RESET_B(net198),
    .D(_0133_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6525_ (.RESET_B(net197),
    .D(net1098),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6526_ (.RESET_B(net196),
    .D(_0135_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _6527_ (.RESET_B(net195),
    .D(net1453),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][3] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _6528_ (.RESET_B(net194),
    .D(net1376),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][4] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6529_ (.RESET_B(net193),
    .D(_0138_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][5] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6530_ (.RESET_B(net192),
    .D(_0139_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][6] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6531_ (.RESET_B(net191),
    .D(_0140_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][7] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6532_ (.RESET_B(net190),
    .D(_0141_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6533_ (.RESET_B(net189),
    .D(_0142_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6534_ (.RESET_B(net188),
    .D(_0143_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[2] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6535_ (.RESET_B(net187),
    .D(net1159),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[3] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6536_ (.RESET_B(net186),
    .D(net1288),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[10] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6537_ (.RESET_B(net185),
    .D(net987),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][0] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6538_ (.RESET_B(net184),
    .D(net997),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6539_ (.RESET_B(net183),
    .D(net1226),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][2] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6540_ (.RESET_B(net182),
    .D(net1207),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][3] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6541_ (.RESET_B(net181),
    .D(_0150_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][4] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6542_ (.RESET_B(net180),
    .D(_0151_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][5] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6543_ (.RESET_B(net179),
    .D(_0152_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][6] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _6544_ (.RESET_B(net178),
    .D(net1333),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][7] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6545_ (.RESET_B(net177),
    .D(_0154_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][8] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6546_ (.RESET_B(net176),
    .D(net1478),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][9] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _6547_ (.RESET_B(net175),
    .D(_0156_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][10] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6548_ (.RESET_B(net174),
    .D(net1170),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][11] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6549_ (.RESET_B(net173),
    .D(net1263),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][12] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6550_ (.RESET_B(net172),
    .D(_0159_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _6551_ (.RESET_B(net171),
    .D(_0160_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6552_ (.RESET_B(net170),
    .D(_0161_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6553_ (.RESET_B(net169),
    .D(_0162_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][3] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6554_ (.RESET_B(net168),
    .D(net1039),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][4] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6555_ (.RESET_B(net167),
    .D(_0164_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][5] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6556_ (.RESET_B(net166),
    .D(_0165_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][6] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6557_ (.RESET_B(net165),
    .D(net1136),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][7] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _6558_ (.RESET_B(net164),
    .D(net1088),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][8] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6559_ (.RESET_B(net163),
    .D(_0168_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][9] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _6560_ (.RESET_B(net162),
    .D(_0169_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][10] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _6561_ (.RESET_B(net161),
    .D(net833),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].z_sign ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _6562_ (.RESET_B(net160),
    .D(_0171_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6563_ (.RESET_B(net159),
    .D(net1166),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6564_ (.RESET_B(net158),
    .D(_0173_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][2] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6565_ (.RESET_B(net157),
    .D(net1353),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][3] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6566_ (.RESET_B(net156),
    .D(net1213),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][4] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6567_ (.RESET_B(net155),
    .D(_0176_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][5] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6568_ (.RESET_B(net154),
    .D(net1254),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][6] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6569_ (.RESET_B(net153),
    .D(net1191),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][7] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6570_ (.RESET_B(net152),
    .D(_0179_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][8] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6571_ (.RESET_B(net151),
    .D(_0180_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6572_ (.RESET_B(net150),
    .D(_0181_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6573_ (.RESET_B(net149),
    .D(net1178),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[2] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _6574_ (.RESET_B(net148),
    .D(net873),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[10] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6575_ (.RESET_B(net147),
    .D(net995),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6576_ (.RESET_B(net146),
    .D(net1018),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _6577_ (.RESET_B(net145),
    .D(net1440),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][2] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6578_ (.RESET_B(net144),
    .D(net1312),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][3] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6579_ (.RESET_B(net143),
    .D(_0188_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][4] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _6580_ (.RESET_B(net142),
    .D(net1294),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][5] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6581_ (.RESET_B(net141),
    .D(_0190_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][6] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6582_ (.RESET_B(net140),
    .D(_0191_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][7] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6583_ (.RESET_B(net139),
    .D(net1460),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][8] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6584_ (.RESET_B(net138),
    .D(_0193_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][9] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6585_ (.RESET_B(net137),
    .D(_0194_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][10] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6586_ (.RESET_B(net136),
    .D(net1274),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][11] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _6587_ (.RESET_B(net135),
    .D(net1400),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][12] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _6588_ (.RESET_B(net134),
    .D(net1143),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].z_sign ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6589_ (.RESET_B(net133),
    .D(_0198_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6590_ (.RESET_B(net132),
    .D(net1366),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6591_ (.RESET_B(net131),
    .D(_0200_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][2] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6592_ (.RESET_B(net130),
    .D(_0201_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][3] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6593_ (.RESET_B(net129),
    .D(_0202_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][4] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6594_ (.RESET_B(net128),
    .D(net1239),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][5] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _6595_ (.RESET_B(net127),
    .D(_0204_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][6] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _6596_ (.RESET_B(net126),
    .D(net1092),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][7] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6597_ (.RESET_B(net125),
    .D(_0206_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][8] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6598_ (.RESET_B(net124),
    .D(_0207_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][9] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6599_ (.RESET_B(net123),
    .D(_0208_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _6600_ (.RESET_B(net122),
    .D(_0209_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _6601_ (.RESET_B(net121),
    .D(net1203),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[10] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6602_ (.RESET_B(net120),
    .D(net1000),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6603_ (.RESET_B(net119),
    .D(net1045),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6604_ (.RESET_B(net118),
    .D(_0213_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][2] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _6605_ (.RESET_B(net117),
    .D(net1448),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][3] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6606_ (.RESET_B(net116),
    .D(_0215_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][4] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6607_ (.RESET_B(net115),
    .D(net1168),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][5] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6608_ (.RESET_B(net114),
    .D(_0217_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][6] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6609_ (.RESET_B(net113),
    .D(net1252),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][7] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6610_ (.RESET_B(net112),
    .D(_0219_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][8] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6611_ (.RESET_B(net111),
    .D(net1174),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][9] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6612_ (.RESET_B(net110),
    .D(_0221_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][10] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6613_ (.RESET_B(net109),
    .D(net1342),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][11] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _6614_ (.RESET_B(net108),
    .D(net1216),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][12] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _6615_ (.RESET_B(net107),
    .D(_0224_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][0] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6616_ (.RESET_B(net106),
    .D(net1161),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6617_ (.RESET_B(net105),
    .D(_0226_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6618_ (.RESET_B(net104),
    .D(net1466),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6619_ (.RESET_B(net103),
    .D(_0228_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][4] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6620_ (.RESET_B(net102),
    .D(net1113),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][5] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6621_ (.RESET_B(net101),
    .D(_0230_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][6] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6622_ (.RESET_B(net100),
    .D(net1123),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][7] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6623_ (.RESET_B(net99),
    .D(_0232_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][8] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6624_ (.RESET_B(net98),
    .D(net1187),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][9] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6625_ (.RESET_B(net97),
    .D(_0234_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][10] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6626_ (.RESET_B(net96),
    .D(_0235_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][11] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6627_ (.RESET_B(net95),
    .D(net990),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6628_ (.RESET_B(net94),
    .D(net1053),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][1] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6629_ (.RESET_B(net93),
    .D(net1490),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6630_ (.RESET_B(net92),
    .D(_0239_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6631_ (.RESET_B(net91),
    .D(_0240_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][4] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6632_ (.RESET_B(net90),
    .D(net1397),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][5] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6633_ (.RESET_B(net89),
    .D(net1561),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][6] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6634_ (.RESET_B(net88),
    .D(net1431),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][7] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _6635_ (.RESET_B(net87),
    .D(net1221),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][8] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _6636_ (.RESET_B(net86),
    .D(_0245_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][9] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6637_ (.RESET_B(net85),
    .D(_0246_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][10] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6638_ (.RESET_B(net84),
    .D(net1198),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][11] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _6639_ (.RESET_B(net83),
    .D(_0248_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt_sum[5] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6640_ (.RESET_B(net82),
    .D(_0249_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6641_ (.RESET_B(net81),
    .D(_0250_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[2] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6642_ (.RESET_B(net80),
    .D(_0251_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[3] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6643_ (.RESET_B(net79),
    .D(_0252_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6644_ (.RESET_B(net78),
    .D(_0253_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[5] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6645_ (.RESET_B(net77),
    .D(_0254_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[6] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6646_ (.RESET_B(net76),
    .D(_0255_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[7] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6647_ (.RESET_B(net75),
    .D(_0256_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[8] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6648_ (.RESET_B(net74),
    .D(_0257_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[9] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6649_ (.RESET_B(net73),
    .D(_0258_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[10] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6650_ (.RESET_B(net72),
    .D(_0259_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[11] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6651_ (.RESET_B(net71),
    .D(_0260_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.freq_reg[12] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _6652_ (.RESET_B(net70),
    .D(_0261_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp[0] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6653_ (.RESET_B(net69),
    .D(net1035),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6654_ (.RESET_B(net68),
    .D(net1102),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][1] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _6655_ (.RESET_B(net67),
    .D(net1395),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][2] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6656_ (.RESET_B(net66),
    .D(_0265_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][3] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6657_ (.RESET_B(net65),
    .D(_0266_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][4] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6658_ (.RESET_B(net64),
    .D(net1276),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][5] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _6659_ (.RESET_B(net63),
    .D(net1164),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][6] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _6660_ (.RESET_B(net62),
    .D(_0269_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][7] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _6661_ (.RESET_B(net61),
    .D(_0270_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][8] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _6662_ (.RESET_B(net60),
    .D(net1290),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][9] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _6663_ (.RESET_B(net59),
    .D(_0272_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][10] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _6664_ (.RESET_B(net58),
    .D(net1292),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][11] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _6665_ (.RESET_B(net57),
    .D(net1409),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][12] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6666_ (.RESET_B(net56),
    .D(_0275_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][0] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6667_ (.RESET_B(net55),
    .D(net1064),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][1] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6668_ (.RESET_B(net54),
    .D(_0277_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][2] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6669_ (.RESET_B(net53),
    .D(net1246),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][3] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6670_ (.RESET_B(net52),
    .D(_0279_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][4] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _6671_ (.RESET_B(net51),
    .D(_0280_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][5] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _6672_ (.RESET_B(net50),
    .D(_0281_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _6673_ (.RESET_B(net49),
    .D(net1540),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[1] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _6674_ (.RESET_B(net48),
    .D(_0283_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[2] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _6675_ (.RESET_B(net47),
    .D(net1182),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[3] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _6676_ (.RESET_B(net46),
    .D(_0285_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[4] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6677_ (.RESET_B(net45),
    .D(net1229),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[5] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _6678_ (.RESET_B(net44),
    .D(net1316),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[10] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _6679_ (.RESET_B(net43),
    .D(_0288_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _6680_ (.RESET_B(net42),
    .D(_0289_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][1] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _6681_ (.RESET_B(net41),
    .D(_0290_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][2] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6682_ (.RESET_B(net40),
    .D(_0291_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][3] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6683_ (.RESET_B(net756),
    .D(net1096),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][4] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _6684_ (.RESET_B(net755),
    .D(_0293_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][5] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _6685_ (.RESET_B(net754),
    .D(net1145),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][6] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6686_ (.RESET_B(net753),
    .D(_0295_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][7] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6687_ (.RESET_B(net752),
    .D(_0296_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][8] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _6688_ (.RESET_B(net751),
    .D(net1270),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][9] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6689_ (.RESET_B(net750),
    .D(_0298_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][10] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _6690_ (.RESET_B(net749),
    .D(net838),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].z_sign ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _6691_ (.RESET_B(net748),
    .D(net972),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6692_ (.RESET_B(net747),
    .D(net1009),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6693_ (.RESET_B(net746),
    .D(net1518),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][2] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6694_ (.RESET_B(net745),
    .D(net1257),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][3] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6695_ (.RESET_B(net744),
    .D(_0304_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][4] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _6696_ (.RESET_B(net743),
    .D(net1418),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][5] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _6697_ (.RESET_B(net742),
    .D(_0306_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][6] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6698_ (.RESET_B(net741),
    .D(net1445),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][7] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _6699_ (.RESET_B(net740),
    .D(_0308_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][8] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _6700_ (.RESET_B(net739),
    .D(net1391),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][9] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _6701_ (.RESET_B(net724),
    .D(_0310_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][10] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _6702_ (.RESET_B(net723),
    .D(net1387),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][11] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _6703_ (.RESET_B(net722),
    .D(net1234),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][12] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6704_ (.RESET_B(net721),
    .D(_0313_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6705_ (.RESET_B(net720),
    .D(net1305),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][1] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6706_ (.RESET_B(net719),
    .D(_0315_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][2] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6707_ (.RESET_B(net718),
    .D(net1368),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][3] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _6708_ (.RESET_B(net717),
    .D(_0317_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][4] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _6709_ (.RESET_B(net716),
    .D(_0318_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[0] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _6710_ (.RESET_B(net715),
    .D(_0319_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _6711_ (.RESET_B(net714),
    .D(net1389),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[2] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _6712_ (.RESET_B(net713),
    .D(_0321_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[3] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _6713_ (.RESET_B(net712),
    .D(net1503),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[4] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _6714_ (.RESET_B(net711),
    .D(_0323_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[5] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _6715_ (.RESET_B(net710),
    .D(_0324_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[6] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6716_ (.RESET_B(net709),
    .D(net1286),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[10] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _6717_ (.RESET_B(net708),
    .D(_0326_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][0] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _6718_ (.RESET_B(net707),
    .D(net853),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _6719_ (.RESET_B(net706),
    .D(net1075),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][2] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _6720_ (.RESET_B(net705),
    .D(_0329_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6721_ (.RESET_B(net704),
    .D(net1090),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][4] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _6722_ (.RESET_B(net703),
    .D(net1359),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][5] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _6723_ (.RESET_B(net702),
    .D(_0332_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][6] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6724_ (.RESET_B(net701),
    .D(net1157),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][7] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _6725_ (.RESET_B(net700),
    .D(_0334_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][8] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _6726_ (.RESET_B(net699),
    .D(_0335_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][9] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _6727_ (.RESET_B(net698),
    .D(net1126),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][10] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6728_ (.RESET_B(net697),
    .D(net812),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].z_sign ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6729_ (.RESET_B(net696),
    .D(net935),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][0] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6730_ (.RESET_B(net695),
    .D(net1232),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6731_ (.RESET_B(net694),
    .D(net1303),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][2] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6732_ (.RESET_B(net693),
    .D(_0341_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][3] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _6733_ (.RESET_B(net692),
    .D(_0342_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][4] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _6734_ (.RESET_B(net691),
    .D(net1416),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][5] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6735_ (.RESET_B(net690),
    .D(net1414),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][6] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _6736_ (.RESET_B(net689),
    .D(net1403),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][7] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6737_ (.RESET_B(net688),
    .D(net1336),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][8] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _6738_ (.RESET_B(net687),
    .D(_0347_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][9] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _6739_ (.RESET_B(net686),
    .D(net1469),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][10] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _6740_ (.RESET_B(net685),
    .D(net1195),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][11] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _6741_ (.RESET_B(net684),
    .D(_0350_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][12] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6742_ (.RESET_B(net683),
    .D(_0351_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[4][0] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6743_ (.RESET_B(net682),
    .D(net1241),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[4][1] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6744_ (.RESET_B(net681),
    .D(_0353_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[4][2] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _6745_ (.RESET_B(net680),
    .D(_0354_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[4][3] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _6746_ (.RESET_B(net679),
    .D(_0355_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[0] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _6747_ (.RESET_B(net678),
    .D(net1378),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[1] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _6748_ (.RESET_B(net677),
    .D(_0357_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[2] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _6749_ (.RESET_B(net676),
    .D(_0358_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[3] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _6750_ (.RESET_B(net675),
    .D(net1521),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[4] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _6751_ (.RESET_B(net674),
    .D(net1451),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[5] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _6752_ (.RESET_B(net673),
    .D(_0361_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[6] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _6753_ (.RESET_B(net672),
    .D(net1119),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[7] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _6754_ (.RESET_B(net671),
    .D(net905),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[10] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _6755_ (.RESET_B(net670),
    .D(_0364_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6756_ (.RESET_B(net669),
    .D(_0365_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6757_ (.RESET_B(net668),
    .D(_0366_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6758_ (.RESET_B(net667),
    .D(_0367_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][3] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _6759_ (.RESET_B(net666),
    .D(net1205),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][4] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6760_ (.RESET_B(net665),
    .D(net1085),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][5] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6761_ (.RESET_B(net664),
    .D(_0370_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][6] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6762_ (.RESET_B(net663),
    .D(net1079),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][7] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6763_ (.RESET_B(net662),
    .D(_0372_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][8] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6764_ (.RESET_B(net661),
    .D(_0373_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][9] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _6765_ (.RESET_B(net660),
    .D(net1129),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][10] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _6766_ (.RESET_B(net659),
    .D(net827),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].z_sign ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _6767_ (.RESET_B(net658),
    .D(net1016),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][0] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6768_ (.RESET_B(net657),
    .D(net1244),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6769_ (.RESET_B(net656),
    .D(net1429),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][2] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _6770_ (.RESET_B(net655),
    .D(net1476),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][3] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _6771_ (.RESET_B(net654),
    .D(net1349),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][4] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6772_ (.RESET_B(net653),
    .D(_0381_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][5] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _6773_ (.RESET_B(net652),
    .D(net1308),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][6] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _6774_ (.RESET_B(net651),
    .D(net1572),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][7] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _6775_ (.RESET_B(net650),
    .D(_0384_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][8] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6776_ (.RESET_B(net649),
    .D(net1328),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][9] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6777_ (.RESET_B(net648),
    .D(net1424),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][10] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _6778_ (.RESET_B(net647),
    .D(_0387_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][11] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6779_ (.RESET_B(net646),
    .D(net1218),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][12] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _6780_ (.RESET_B(net645),
    .D(_0389_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[3][0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6781_ (.RESET_B(net644),
    .D(net1148),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[3][1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6782_ (.RESET_B(net643),
    .D(_0391_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[3][2] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _6783_ (.RESET_B(net642),
    .D(net1511),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _6784_ (.RESET_B(net641),
    .D(net1250),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _6785_ (.RESET_B(net640),
    .D(_0394_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[2] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _6786_ (.RESET_B(net639),
    .D(_0395_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[3] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6787_ (.RESET_B(net638),
    .D(net1555),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[4] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6788_ (.RESET_B(net637),
    .D(net1437),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[5] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6789_ (.RESET_B(net636),
    .D(_0398_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[6] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6790_ (.RESET_B(net635),
    .D(_0399_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[7] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _6791_ (.RESET_B(net634),
    .D(_0400_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[8] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _6792_ (.RESET_B(net633),
    .D(net1324),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[10] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6793_ (.RESET_B(net632),
    .D(_0402_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6794_ (.RESET_B(net631),
    .D(_0403_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6795_ (.RESET_B(net630),
    .D(_0404_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6796_ (.RESET_B(net629),
    .D(_0405_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _6797_ (.RESET_B(net628),
    .D(_0406_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][4] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6798_ (.RESET_B(net627),
    .D(_0407_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][5] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6799_ (.RESET_B(net626),
    .D(_0408_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6800_ (.RESET_B(net625),
    .D(_0409_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][7] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6801_ (.RESET_B(net624),
    .D(_0410_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][8] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6802_ (.RESET_B(net623),
    .D(net1155),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][9] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6803_ (.RESET_B(net622),
    .D(_0412_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][10] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _6804_ (.RESET_B(net621),
    .D(_0413_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].z_sign ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6805_ (.RESET_B(net620),
    .D(net1048),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6806_ (.RESET_B(net619),
    .D(net1077),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _6807_ (.RESET_B(net618),
    .D(_0416_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][2] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _6808_ (.RESET_B(net617),
    .D(net1340),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][3] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _6809_ (.RESET_B(net616),
    .D(net1297),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][4] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6810_ (.RESET_B(net615),
    .D(net1211),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][5] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _6811_ (.RESET_B(net614),
    .D(_0420_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][6] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _6812_ (.RESET_B(net613),
    .D(_0421_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][7] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _6813_ (.RESET_B(net612),
    .D(net1321),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][8] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _6814_ (.RESET_B(net611),
    .D(_0423_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][9] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _6815_ (.RESET_B(net610),
    .D(net1373),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6816_ (.RESET_B(net609),
    .D(_0425_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][11] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6817_ (.RESET_B(net608),
    .D(net1132),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][12] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6818_ (.RESET_B(net607),
    .D(_0427_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[2][0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _6819_ (.RESET_B(net606),
    .D(_0428_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[2][1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _6820_ (.RESET_B(net605),
    .D(_0429_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[0] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _6821_ (.RESET_B(net604),
    .D(net1299),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[1] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _6822_ (.RESET_B(net603),
    .D(_0431_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[2] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _6823_ (.RESET_B(net602),
    .D(net1407),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[3] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_2 _6824_ (.RESET_B(net601),
    .D(_0433_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[4] ),
    .CLK(clknet_leaf_60_clk));
 sg13g2_dfrbpq_1 _6825_ (.RESET_B(net600),
    .D(_0434_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[5] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _6826_ (.RESET_B(net599),
    .D(_0435_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[6] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _6827_ (.RESET_B(net598),
    .D(net1492),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[7] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _6828_ (.RESET_B(net597),
    .D(_0437_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[8] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6829_ (.RESET_B(net596),
    .D(net1345),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[9] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6830_ (.RESET_B(net595),
    .D(net1283),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[10] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6831_ (.RESET_B(net594),
    .D(net762),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6832_ (.RESET_B(net593),
    .D(_0441_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _6833_ (.RESET_B(net592),
    .D(_0442_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][2] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6834_ (.RESET_B(net591),
    .D(_0443_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6835_ (.RESET_B(net590),
    .D(net1050),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][4] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6836_ (.RESET_B(net589),
    .D(net1331),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][5] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6837_ (.RESET_B(net588),
    .D(net1236),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][6] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _6838_ (.RESET_B(net587),
    .D(_0447_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][7] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6839_ (.RESET_B(net586),
    .D(_0448_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][8] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6840_ (.RESET_B(net585),
    .D(net1073),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][9] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6841_ (.RESET_B(net584),
    .D(_0450_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][10] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _6842_ (.RESET_B(net583),
    .D(_0451_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].z_sign ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _6843_ (.RESET_B(net582),
    .D(net969),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _6844_ (.RESET_B(net581),
    .D(_0453_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][1] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _6845_ (.RESET_B(net580),
    .D(_0454_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][2] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _6846_ (.RESET_B(net579),
    .D(_0455_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][3] ),
    .CLK(clknet_leaf_65_clk));
 sg13g2_dfrbpq_2 _6847_ (.RESET_B(net578),
    .D(_0456_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][4] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _6848_ (.RESET_B(net577),
    .D(_0457_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][5] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _6849_ (.RESET_B(net576),
    .D(_0458_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][6] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _6850_ (.RESET_B(net575),
    .D(_0459_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][7] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _6851_ (.RESET_B(net570),
    .D(_0460_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][8] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _6852_ (.RESET_B(net568),
    .D(_0461_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][9] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6853_ (.RESET_B(net566),
    .D(_0462_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][10] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _6854_ (.RESET_B(net562),
    .D(_0463_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][11] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6855_ (.RESET_B(net560),
    .D(_0464_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][12] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6856_ (.RESET_B(net557),
    .D(_0465_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[0] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _6857_ (.RESET_B(net371),
    .D(_0466_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[1] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _6858_ (.RESET_B(net369),
    .D(_0467_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[2] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_1 _6859_ (.RESET_B(net367),
    .D(_0468_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[3] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _6860_ (.RESET_B(net365),
    .D(net1042),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[4] ),
    .CLK(clknet_leaf_64_clk));
 sg13g2_dfrbpq_2 _6861_ (.RESET_B(net363),
    .D(_0470_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[5] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _6862_ (.RESET_B(net361),
    .D(_0471_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[6] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _6863_ (.RESET_B(net359),
    .D(_0472_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[7] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _6864_ (.RESET_B(net357),
    .D(_0473_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[8] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6865_ (.RESET_B(net355),
    .D(_0474_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[9] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6866_ (.RESET_B(net353),
    .D(_0475_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _6867_ (.RESET_B(net351),
    .D(_0476_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[11] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _6868_ (.RESET_B(net349),
    .D(_0477_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6869_ (.RESET_B(net347),
    .D(_0478_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6870_ (.RESET_B(net345),
    .D(_0479_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][2] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6871_ (.RESET_B(net343),
    .D(_0480_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6872_ (.RESET_B(net341),
    .D(_0481_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][4] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6873_ (.RESET_B(net339),
    .D(_0482_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][5] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6874_ (.RESET_B(net337),
    .D(_0483_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][6] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6875_ (.RESET_B(net335),
    .D(_0484_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][7] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _6876_ (.RESET_B(net333),
    .D(_0485_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][8] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _6877_ (.RESET_B(net331),
    .D(_0486_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][9] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6878_ (.RESET_B(net329),
    .D(_0487_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][10] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6879_ (.RESET_B(net327),
    .D(net816),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].z_sign ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _6880_ (.RESET_B(net325),
    .D(_0489_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[0] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6881_ (.RESET_B(net323),
    .D(_0490_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6882_ (.RESET_B(net321),
    .D(_0491_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[2] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6883_ (.RESET_B(net319),
    .D(_0492_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _6884_ (.RESET_B(net317),
    .D(_0493_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[4] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _6885_ (.RESET_B(net315),
    .D(_0494_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[5] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6886_ (.RESET_B(net300),
    .D(_0495_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[6] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _6887_ (.RESET_B(net298),
    .D(net797),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[7] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6888_ (.RESET_B(net296),
    .D(_0497_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6889_ (.RESET_B(net294),
    .D(_0498_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[9] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6890_ (.RESET_B(net292),
    .D(_0499_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[10] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _6891_ (.RESET_B(net726),
    .D(_0500_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.SINout[11] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _6892_ (.RESET_B(net727),
    .D(net442),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.x_start[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _6893_ (.RESET_B(net728),
    .D(_0519_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][0] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6894_ (.RESET_B(net729),
    .D(_0522_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6895_ (.RESET_B(net730),
    .D(_0523_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][2] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _6896_ (.RESET_B(net731),
    .D(net850),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6897_ (.RESET_B(net732),
    .D(_0525_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][4] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _6898_ (.RESET_B(net733),
    .D(_0526_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][5] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _6899_ (.RESET_B(net734),
    .D(_0527_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][6] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6900_ (.RESET_B(net735),
    .D(_0528_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6901_ (.RESET_B(net736),
    .D(_0529_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][8] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _6902_ (.RESET_B(net737),
    .D(_0530_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][9] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _6903_ (.RESET_B(net738),
    .D(_0520_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][10] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _6904_ (.RESET_B(net250),
    .D(_0521_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[0].z_sign ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _6905_ (.RESET_B(net290),
    .D(net1),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.resetn ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _6906_ (.RESET_B(net288),
    .D(_0501_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6907_ (.RESET_B(net286),
    .D(_0502_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6908_ (.RESET_B(net284),
    .D(net900),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6909_ (.RESET_B(net282),
    .D(_0504_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[3] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _6910_ (.RESET_B(net280),
    .D(net928),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[4] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _6911_ (.RESET_B(net278),
    .D(net845),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[5] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6912_ (.RESET_B(net276),
    .D(_0507_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[6] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6913_ (.RESET_B(net272),
    .D(net1109),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _6914_ (.RESET_B(net270),
    .D(_0509_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[8] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _6915_ (.RESET_B(net268),
    .D(net848),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[9] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6916_ (.RESET_B(net266),
    .D(_0511_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[10] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6917_ (.RESET_B(net264),
    .D(_0512_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[11] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6918_ (.RESET_B(net262),
    .D(_0513_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[12] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _6919_ (.RESET_B(net260),
    .D(net960),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[13] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _6920_ (.RESET_B(net258),
    .D(_0515_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[14] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6921_ (.RESET_B(net256),
    .D(net855),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[15] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _6922_ (.RESET_B(net254),
    .D(_0517_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[16] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _6923_ (.RESET_B(net252),
    .D(_0518_),
    .Q(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[17] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_tiehi _6681__41 (.L_HI(net41));
 sg13g2_tiehi _6680__42 (.L_HI(net42));
 sg13g2_tiehi _6679__43 (.L_HI(net43));
 sg13g2_tiehi _6678__44 (.L_HI(net44));
 sg13g2_tiehi _6677__45 (.L_HI(net45));
 sg13g2_tiehi _6676__46 (.L_HI(net46));
 sg13g2_tiehi _6675__47 (.L_HI(net47));
 sg13g2_tiehi _6674__48 (.L_HI(net48));
 sg13g2_tiehi _6673__49 (.L_HI(net49));
 sg13g2_tiehi _6672__50 (.L_HI(net50));
 sg13g2_tiehi _6671__51 (.L_HI(net51));
 sg13g2_tiehi _6670__52 (.L_HI(net52));
 sg13g2_tiehi _6669__53 (.L_HI(net53));
 sg13g2_tiehi _6668__54 (.L_HI(net54));
 sg13g2_tiehi _6667__55 (.L_HI(net55));
 sg13g2_tiehi _6666__56 (.L_HI(net56));
 sg13g2_tiehi _6665__57 (.L_HI(net57));
 sg13g2_tiehi _6664__58 (.L_HI(net58));
 sg13g2_tiehi _6663__59 (.L_HI(net59));
 sg13g2_tiehi _6662__60 (.L_HI(net60));
 sg13g2_tiehi _6661__61 (.L_HI(net61));
 sg13g2_tiehi _6660__62 (.L_HI(net62));
 sg13g2_tiehi _6659__63 (.L_HI(net63));
 sg13g2_tiehi _6658__64 (.L_HI(net64));
 sg13g2_tiehi _6657__65 (.L_HI(net65));
 sg13g2_tiehi _6656__66 (.L_HI(net66));
 sg13g2_tiehi _6655__67 (.L_HI(net67));
 sg13g2_tiehi _6654__68 (.L_HI(net68));
 sg13g2_tiehi _6653__69 (.L_HI(net69));
 sg13g2_tiehi _6652__70 (.L_HI(net70));
 sg13g2_tiehi _6651__71 (.L_HI(net71));
 sg13g2_tiehi _6650__72 (.L_HI(net72));
 sg13g2_tiehi _6649__73 (.L_HI(net73));
 sg13g2_tiehi _6648__74 (.L_HI(net74));
 sg13g2_tiehi _6647__75 (.L_HI(net75));
 sg13g2_tiehi _6646__76 (.L_HI(net76));
 sg13g2_tiehi _6645__77 (.L_HI(net77));
 sg13g2_tiehi _6644__78 (.L_HI(net78));
 sg13g2_tiehi _6643__79 (.L_HI(net79));
 sg13g2_tiehi _6642__80 (.L_HI(net80));
 sg13g2_tiehi _6641__81 (.L_HI(net81));
 sg13g2_tiehi _6640__82 (.L_HI(net82));
 sg13g2_tiehi _6639__83 (.L_HI(net83));
 sg13g2_tiehi _6638__84 (.L_HI(net84));
 sg13g2_tiehi _6637__85 (.L_HI(net85));
 sg13g2_tiehi _6636__86 (.L_HI(net86));
 sg13g2_tiehi _6635__87 (.L_HI(net87));
 sg13g2_tiehi _6634__88 (.L_HI(net88));
 sg13g2_tiehi _6633__89 (.L_HI(net89));
 sg13g2_tiehi _6632__90 (.L_HI(net90));
 sg13g2_tiehi _6631__91 (.L_HI(net91));
 sg13g2_tiehi _6630__92 (.L_HI(net92));
 sg13g2_tiehi _6629__93 (.L_HI(net93));
 sg13g2_tiehi _6628__94 (.L_HI(net94));
 sg13g2_tiehi _6627__95 (.L_HI(net95));
 sg13g2_tiehi _6626__96 (.L_HI(net96));
 sg13g2_tiehi _6625__97 (.L_HI(net97));
 sg13g2_tiehi _6624__98 (.L_HI(net98));
 sg13g2_tiehi _6623__99 (.L_HI(net99));
 sg13g2_tiehi _6622__100 (.L_HI(net100));
 sg13g2_tiehi _6621__101 (.L_HI(net101));
 sg13g2_tiehi _6620__102 (.L_HI(net102));
 sg13g2_tiehi _6619__103 (.L_HI(net103));
 sg13g2_tiehi _6618__104 (.L_HI(net104));
 sg13g2_tiehi _6617__105 (.L_HI(net105));
 sg13g2_tiehi _6616__106 (.L_HI(net106));
 sg13g2_tiehi _6615__107 (.L_HI(net107));
 sg13g2_tiehi _6614__108 (.L_HI(net108));
 sg13g2_tiehi _6613__109 (.L_HI(net109));
 sg13g2_tiehi _6612__110 (.L_HI(net110));
 sg13g2_tiehi _6611__111 (.L_HI(net111));
 sg13g2_tiehi _6610__112 (.L_HI(net112));
 sg13g2_tiehi _6609__113 (.L_HI(net113));
 sg13g2_tiehi _6608__114 (.L_HI(net114));
 sg13g2_tiehi _6607__115 (.L_HI(net115));
 sg13g2_tiehi _6606__116 (.L_HI(net116));
 sg13g2_tiehi _6605__117 (.L_HI(net117));
 sg13g2_tiehi _6604__118 (.L_HI(net118));
 sg13g2_tiehi _6603__119 (.L_HI(net119));
 sg13g2_tiehi _6602__120 (.L_HI(net120));
 sg13g2_tiehi _6601__121 (.L_HI(net121));
 sg13g2_tiehi _6600__122 (.L_HI(net122));
 sg13g2_tiehi _6599__123 (.L_HI(net123));
 sg13g2_tiehi _6598__124 (.L_HI(net124));
 sg13g2_tiehi _6597__125 (.L_HI(net125));
 sg13g2_tiehi _6596__126 (.L_HI(net126));
 sg13g2_tiehi _6595__127 (.L_HI(net127));
 sg13g2_tiehi _6594__128 (.L_HI(net128));
 sg13g2_tiehi _6593__129 (.L_HI(net129));
 sg13g2_tiehi _6592__130 (.L_HI(net130));
 sg13g2_tiehi _6591__131 (.L_HI(net131));
 sg13g2_tiehi _6590__132 (.L_HI(net132));
 sg13g2_tiehi _6589__133 (.L_HI(net133));
 sg13g2_tiehi _6588__134 (.L_HI(net134));
 sg13g2_tiehi _6587__135 (.L_HI(net135));
 sg13g2_tiehi _6586__136 (.L_HI(net136));
 sg13g2_tiehi _6585__137 (.L_HI(net137));
 sg13g2_tiehi _6584__138 (.L_HI(net138));
 sg13g2_tiehi _6583__139 (.L_HI(net139));
 sg13g2_tiehi _6582__140 (.L_HI(net140));
 sg13g2_tiehi _6581__141 (.L_HI(net141));
 sg13g2_tiehi _6580__142 (.L_HI(net142));
 sg13g2_tiehi _6579__143 (.L_HI(net143));
 sg13g2_tiehi _6578__144 (.L_HI(net144));
 sg13g2_tiehi _6577__145 (.L_HI(net145));
 sg13g2_tiehi _6576__146 (.L_HI(net146));
 sg13g2_tiehi _6575__147 (.L_HI(net147));
 sg13g2_tiehi _6574__148 (.L_HI(net148));
 sg13g2_tiehi _6573__149 (.L_HI(net149));
 sg13g2_tiehi _6572__150 (.L_HI(net150));
 sg13g2_tiehi _6571__151 (.L_HI(net151));
 sg13g2_tiehi _6570__152 (.L_HI(net152));
 sg13g2_tiehi _6569__153 (.L_HI(net153));
 sg13g2_tiehi _6568__154 (.L_HI(net154));
 sg13g2_tiehi _6567__155 (.L_HI(net155));
 sg13g2_tiehi _6566__156 (.L_HI(net156));
 sg13g2_tiehi _6565__157 (.L_HI(net157));
 sg13g2_tiehi _6564__158 (.L_HI(net158));
 sg13g2_tiehi _6563__159 (.L_HI(net159));
 sg13g2_tiehi _6562__160 (.L_HI(net160));
 sg13g2_tiehi _6561__161 (.L_HI(net161));
 sg13g2_tiehi _6560__162 (.L_HI(net162));
 sg13g2_tiehi _6559__163 (.L_HI(net163));
 sg13g2_tiehi _6558__164 (.L_HI(net164));
 sg13g2_tiehi _6557__165 (.L_HI(net165));
 sg13g2_tiehi _6556__166 (.L_HI(net166));
 sg13g2_tiehi _6555__167 (.L_HI(net167));
 sg13g2_tiehi _6554__168 (.L_HI(net168));
 sg13g2_tiehi _6553__169 (.L_HI(net169));
 sg13g2_tiehi _6552__170 (.L_HI(net170));
 sg13g2_tiehi _6551__171 (.L_HI(net171));
 sg13g2_tiehi _6550__172 (.L_HI(net172));
 sg13g2_tiehi _6549__173 (.L_HI(net173));
 sg13g2_tiehi _6548__174 (.L_HI(net174));
 sg13g2_tiehi _6547__175 (.L_HI(net175));
 sg13g2_tiehi _6546__176 (.L_HI(net176));
 sg13g2_tiehi _6545__177 (.L_HI(net177));
 sg13g2_tiehi _6544__178 (.L_HI(net178));
 sg13g2_tiehi _6543__179 (.L_HI(net179));
 sg13g2_tiehi _6542__180 (.L_HI(net180));
 sg13g2_tiehi _6541__181 (.L_HI(net181));
 sg13g2_tiehi _6540__182 (.L_HI(net182));
 sg13g2_tiehi _6539__183 (.L_HI(net183));
 sg13g2_tiehi _6538__184 (.L_HI(net184));
 sg13g2_tiehi _6537__185 (.L_HI(net185));
 sg13g2_tiehi _6536__186 (.L_HI(net186));
 sg13g2_tiehi _6535__187 (.L_HI(net187));
 sg13g2_tiehi _6534__188 (.L_HI(net188));
 sg13g2_tiehi _6533__189 (.L_HI(net189));
 sg13g2_tiehi _6532__190 (.L_HI(net190));
 sg13g2_tiehi _6531__191 (.L_HI(net191));
 sg13g2_tiehi _6530__192 (.L_HI(net192));
 sg13g2_tiehi _6529__193 (.L_HI(net193));
 sg13g2_tiehi _6528__194 (.L_HI(net194));
 sg13g2_tiehi _6527__195 (.L_HI(net195));
 sg13g2_tiehi _6526__196 (.L_HI(net196));
 sg13g2_tiehi _6525__197 (.L_HI(net197));
 sg13g2_tiehi _6524__198 (.L_HI(net198));
 sg13g2_tiehi _6523__199 (.L_HI(net199));
 sg13g2_tiehi _6522__200 (.L_HI(net200));
 sg13g2_tiehi _6521__201 (.L_HI(net201));
 sg13g2_tiehi _6520__202 (.L_HI(net202));
 sg13g2_tiehi _6519__203 (.L_HI(net203));
 sg13g2_tiehi _6518__204 (.L_HI(net204));
 sg13g2_tiehi _6517__205 (.L_HI(net205));
 sg13g2_tiehi _6516__206 (.L_HI(net206));
 sg13g2_tiehi _6515__207 (.L_HI(net207));
 sg13g2_tiehi _6514__208 (.L_HI(net208));
 sg13g2_tiehi _6513__209 (.L_HI(net209));
 sg13g2_tiehi _6512__210 (.L_HI(net210));
 sg13g2_tiehi _6511__211 (.L_HI(net211));
 sg13g2_tiehi _6510__212 (.L_HI(net212));
 sg13g2_tiehi _6509__213 (.L_HI(net213));
 sg13g2_tiehi _6508__214 (.L_HI(net214));
 sg13g2_tiehi _6507__215 (.L_HI(net215));
 sg13g2_tiehi _6506__216 (.L_HI(net216));
 sg13g2_tiehi _6505__217 (.L_HI(net217));
 sg13g2_tiehi _6504__218 (.L_HI(net218));
 sg13g2_tiehi _6503__219 (.L_HI(net219));
 sg13g2_tiehi _6502__220 (.L_HI(net220));
 sg13g2_tiehi _6501__221 (.L_HI(net221));
 sg13g2_tiehi _6500__222 (.L_HI(net222));
 sg13g2_tiehi _6499__223 (.L_HI(net223));
 sg13g2_tiehi _6498__224 (.L_HI(net224));
 sg13g2_tiehi _6497__225 (.L_HI(net225));
 sg13g2_tiehi _6496__226 (.L_HI(net226));
 sg13g2_tiehi _6495__227 (.L_HI(net227));
 sg13g2_tiehi _6494__228 (.L_HI(net228));
 sg13g2_tiehi _6493__229 (.L_HI(net229));
 sg13g2_tiehi _6492__230 (.L_HI(net230));
 sg13g2_tiehi _6491__231 (.L_HI(net231));
 sg13g2_tiehi _6490__232 (.L_HI(net232));
 sg13g2_tiehi _6489__233 (.L_HI(net233));
 sg13g2_tiehi _6488__234 (.L_HI(net234));
 sg13g2_tiehi _6487__235 (.L_HI(net235));
 sg13g2_tiehi _6486__236 (.L_HI(net236));
 sg13g2_tiehi _6485__237 (.L_HI(net237));
 sg13g2_tiehi _6484__238 (.L_HI(net238));
 sg13g2_tiehi _6483__239 (.L_HI(net239));
 sg13g2_tiehi _6482__240 (.L_HI(net240));
 sg13g2_tiehi _6481__241 (.L_HI(net241));
 sg13g2_tiehi _6480__242 (.L_HI(net242));
 sg13g2_tiehi _6479__243 (.L_HI(net243));
 sg13g2_tiehi _6478__244 (.L_HI(net244));
 sg13g2_tiehi _6477__245 (.L_HI(net245));
 sg13g2_tiehi _6476__246 (.L_HI(net246));
 sg13g2_tiehi _6475__247 (.L_HI(net247));
 sg13g2_tiehi _6474__248 (.L_HI(net248));
 sg13g2_tiehi _6473__249 (.L_HI(net249));
 sg13g2_tiehi _6904__250 (.L_HI(net250));
 sg13g2_tiehi _6472__251 (.L_HI(net251));
 sg13g2_tiehi _6923__252 (.L_HI(net252));
 sg13g2_tiehi _6471__253 (.L_HI(net253));
 sg13g2_tiehi _6922__254 (.L_HI(net254));
 sg13g2_tiehi _6470__255 (.L_HI(net255));
 sg13g2_tiehi _6921__256 (.L_HI(net256));
 sg13g2_tiehi _6469__257 (.L_HI(net257));
 sg13g2_tiehi _6920__258 (.L_HI(net258));
 sg13g2_tiehi _6468__259 (.L_HI(net259));
 sg13g2_tiehi _6919__260 (.L_HI(net260));
 sg13g2_tiehi _6467__261 (.L_HI(net261));
 sg13g2_tiehi _6918__262 (.L_HI(net262));
 sg13g2_tiehi _6466__263 (.L_HI(net263));
 sg13g2_tiehi _6917__264 (.L_HI(net264));
 sg13g2_tiehi _6465__265 (.L_HI(net265));
 sg13g2_tiehi _6916__266 (.L_HI(net266));
 sg13g2_tiehi _6464__267 (.L_HI(net267));
 sg13g2_tiehi _6915__268 (.L_HI(net268));
 sg13g2_tiehi _6463__269 (.L_HI(net269));
 sg13g2_tiehi _6914__270 (.L_HI(net270));
 sg13g2_tiehi _6462__271 (.L_HI(net271));
 sg13g2_tiehi _6913__272 (.L_HI(net272));
 sg13g2_tiehi _6461__273 (.L_HI(net273));
 sg13g2_tiehi _6460__274 (.L_HI(net274));
 sg13g2_tiehi _6459__275 (.L_HI(net275));
 sg13g2_tiehi _6912__276 (.L_HI(net276));
 sg13g2_tiehi _6458__277 (.L_HI(net277));
 sg13g2_tiehi _6911__278 (.L_HI(net278));
 sg13g2_tiehi _6457__279 (.L_HI(net279));
 sg13g2_tiehi _6910__280 (.L_HI(net280));
 sg13g2_tiehi _6456__281 (.L_HI(net281));
 sg13g2_tiehi _6909__282 (.L_HI(net282));
 sg13g2_tiehi _6455__283 (.L_HI(net283));
 sg13g2_tiehi _6908__284 (.L_HI(net284));
 sg13g2_tiehi _6454__285 (.L_HI(net285));
 sg13g2_tiehi _6907__286 (.L_HI(net286));
 sg13g2_tiehi _6453__287 (.L_HI(net287));
 sg13g2_tiehi _6906__288 (.L_HI(net288));
 sg13g2_tiehi _6452__289 (.L_HI(net289));
 sg13g2_tiehi _6905__290 (.L_HI(net290));
 sg13g2_tiehi _6451__291 (.L_HI(net291));
 sg13g2_tiehi _6890__292 (.L_HI(net292));
 sg13g2_tiehi _6450__293 (.L_HI(net293));
 sg13g2_tiehi _6889__294 (.L_HI(net294));
 sg13g2_tiehi _6449__295 (.L_HI(net295));
 sg13g2_tiehi _6888__296 (.L_HI(net296));
 sg13g2_tiehi _6448__297 (.L_HI(net297));
 sg13g2_tiehi _6887__298 (.L_HI(net298));
 sg13g2_tiehi _6447__299 (.L_HI(net299));
 sg13g2_tiehi _6886__300 (.L_HI(net300));
 sg13g2_tiehi _6446__301 (.L_HI(net301));
 sg13g2_tiehi _6445__302 (.L_HI(net302));
 sg13g2_tiehi _6444__303 (.L_HI(net303));
 sg13g2_tiehi _6443__304 (.L_HI(net304));
 sg13g2_tiehi _6442__305 (.L_HI(net305));
 sg13g2_tiehi _6441__306 (.L_HI(net306));
 sg13g2_tiehi _6440__307 (.L_HI(net307));
 sg13g2_tiehi _6439__308 (.L_HI(net308));
 sg13g2_tiehi _6438__309 (.L_HI(net309));
 sg13g2_tiehi _6437__310 (.L_HI(net310));
 sg13g2_tiehi _6436__311 (.L_HI(net311));
 sg13g2_tiehi _6435__312 (.L_HI(net312));
 sg13g2_tiehi _6434__313 (.L_HI(net313));
 sg13g2_tiehi _6433__314 (.L_HI(net314));
 sg13g2_tiehi _6885__315 (.L_HI(net315));
 sg13g2_tiehi _6432__316 (.L_HI(net316));
 sg13g2_tiehi _6884__317 (.L_HI(net317));
 sg13g2_tiehi _6431__318 (.L_HI(net318));
 sg13g2_tiehi _6883__319 (.L_HI(net319));
 sg13g2_tiehi _6430__320 (.L_HI(net320));
 sg13g2_tiehi _6882__321 (.L_HI(net321));
 sg13g2_tiehi _6429__322 (.L_HI(net322));
 sg13g2_tiehi _6881__323 (.L_HI(net323));
 sg13g2_tiehi _6428__324 (.L_HI(net324));
 sg13g2_tiehi _6880__325 (.L_HI(net325));
 sg13g2_tiehi _6427__326 (.L_HI(net326));
 sg13g2_tiehi _6879__327 (.L_HI(net327));
 sg13g2_tiehi _6426__328 (.L_HI(net328));
 sg13g2_tiehi _6878__329 (.L_HI(net329));
 sg13g2_tiehi _6425__330 (.L_HI(net330));
 sg13g2_tiehi _6877__331 (.L_HI(net331));
 sg13g2_tiehi _6424__332 (.L_HI(net332));
 sg13g2_tiehi _6876__333 (.L_HI(net333));
 sg13g2_tiehi _6423__334 (.L_HI(net334));
 sg13g2_tiehi _6875__335 (.L_HI(net335));
 sg13g2_tiehi _6422__336 (.L_HI(net336));
 sg13g2_tiehi _6874__337 (.L_HI(net337));
 sg13g2_tiehi _6421__338 (.L_HI(net338));
 sg13g2_tiehi _6873__339 (.L_HI(net339));
 sg13g2_tiehi _6420__340 (.L_HI(net340));
 sg13g2_tiehi _6872__341 (.L_HI(net341));
 sg13g2_tiehi _6419__342 (.L_HI(net342));
 sg13g2_tiehi _6871__343 (.L_HI(net343));
 sg13g2_tiehi _6418__344 (.L_HI(net344));
 sg13g2_tiehi _6870__345 (.L_HI(net345));
 sg13g2_tiehi _6417__346 (.L_HI(net346));
 sg13g2_tiehi _6869__347 (.L_HI(net347));
 sg13g2_tiehi _6416__348 (.L_HI(net348));
 sg13g2_tiehi _6868__349 (.L_HI(net349));
 sg13g2_tiehi _6415__350 (.L_HI(net350));
 sg13g2_tiehi _6867__351 (.L_HI(net351));
 sg13g2_tiehi _6414__352 (.L_HI(net352));
 sg13g2_tiehi _6866__353 (.L_HI(net353));
 sg13g2_tiehi _6413__354 (.L_HI(net354));
 sg13g2_tiehi _6865__355 (.L_HI(net355));
 sg13g2_tiehi _6412__356 (.L_HI(net356));
 sg13g2_tiehi _6864__357 (.L_HI(net357));
 sg13g2_tiehi _6411__358 (.L_HI(net358));
 sg13g2_tiehi _6863__359 (.L_HI(net359));
 sg13g2_tiehi _6410__360 (.L_HI(net360));
 sg13g2_tiehi _6862__361 (.L_HI(net361));
 sg13g2_tiehi _6409__362 (.L_HI(net362));
 sg13g2_tiehi _6861__363 (.L_HI(net363));
 sg13g2_tiehi _6408__364 (.L_HI(net364));
 sg13g2_tiehi _6860__365 (.L_HI(net365));
 sg13g2_tiehi _6407__366 (.L_HI(net366));
 sg13g2_tiehi _6859__367 (.L_HI(net367));
 sg13g2_tiehi _6406__368 (.L_HI(net368));
 sg13g2_tiehi _6858__369 (.L_HI(net369));
 sg13g2_tiehi _6405__370 (.L_HI(net370));
 sg13g2_tiehi _6857__371 (.L_HI(net371));
 sg13g2_tiehi _6404__372 (.L_HI(net556));
 sg13g2_tiehi _6856__373 (.L_HI(net557));
 sg13g2_tiehi _6403__374 (.L_HI(net558));
 sg13g2_tiehi _6402__375 (.L_HI(net559));
 sg13g2_tiehi _6855__376 (.L_HI(net560));
 sg13g2_tiehi _6401__377 (.L_HI(net561));
 sg13g2_tiehi _6854__378 (.L_HI(net562));
 sg13g2_tiehi _6400__379 (.L_HI(net563));
 sg13g2_tiehi _6399__380 (.L_HI(net564));
 sg13g2_tiehi _6398__381 (.L_HI(net565));
 sg13g2_tiehi _6853__382 (.L_HI(net566));
 sg13g2_tiehi _6397__383 (.L_HI(net567));
 sg13g2_tiehi _6852__384 (.L_HI(net568));
 sg13g2_tiehi _6396__385 (.L_HI(net569));
 sg13g2_tiehi _6851__386 (.L_HI(net570));
 sg13g2_tiehi _6395__387 (.L_HI(net571));
 sg13g2_tiehi _6394__388 (.L_HI(net572));
 sg13g2_tiehi _6393__389 (.L_HI(net573));
 sg13g2_tiehi _6392__390 (.L_HI(net574));
 sg13g2_tiehi _6850__391 (.L_HI(net575));
 sg13g2_tiehi _6849__392 (.L_HI(net576));
 sg13g2_tiehi _6848__393 (.L_HI(net577));
 sg13g2_tiehi _6847__394 (.L_HI(net578));
 sg13g2_tiehi _6846__395 (.L_HI(net579));
 sg13g2_tiehi _6845__396 (.L_HI(net580));
 sg13g2_tiehi _6844__397 (.L_HI(net581));
 sg13g2_tiehi _6843__398 (.L_HI(net582));
 sg13g2_tiehi _6842__399 (.L_HI(net583));
 sg13g2_tiehi _6841__400 (.L_HI(net584));
 sg13g2_tiehi _6840__401 (.L_HI(net585));
 sg13g2_tiehi _6839__402 (.L_HI(net586));
 sg13g2_tiehi _6838__403 (.L_HI(net587));
 sg13g2_tiehi _6837__404 (.L_HI(net588));
 sg13g2_tiehi _6836__405 (.L_HI(net589));
 sg13g2_tiehi _6835__406 (.L_HI(net590));
 sg13g2_tiehi _6834__407 (.L_HI(net591));
 sg13g2_tiehi _6833__408 (.L_HI(net592));
 sg13g2_tiehi _6832__409 (.L_HI(net593));
 sg13g2_tiehi _6831__410 (.L_HI(net594));
 sg13g2_tiehi _6830__411 (.L_HI(net595));
 sg13g2_tiehi _6829__412 (.L_HI(net596));
 sg13g2_tiehi _6828__413 (.L_HI(net597));
 sg13g2_tiehi _6827__414 (.L_HI(net598));
 sg13g2_tiehi _6826__415 (.L_HI(net599));
 sg13g2_tiehi _6825__416 (.L_HI(net600));
 sg13g2_tiehi _6824__417 (.L_HI(net601));
 sg13g2_tiehi _6823__418 (.L_HI(net602));
 sg13g2_tiehi _6822__419 (.L_HI(net603));
 sg13g2_tiehi _6821__420 (.L_HI(net604));
 sg13g2_tiehi _6820__421 (.L_HI(net605));
 sg13g2_tiehi _6819__422 (.L_HI(net606));
 sg13g2_tiehi _6818__423 (.L_HI(net607));
 sg13g2_tiehi _6817__424 (.L_HI(net608));
 sg13g2_tiehi _6816__425 (.L_HI(net609));
 sg13g2_tiehi _6815__426 (.L_HI(net610));
 sg13g2_tiehi _6814__427 (.L_HI(net611));
 sg13g2_tiehi _6813__428 (.L_HI(net612));
 sg13g2_tiehi _6812__429 (.L_HI(net613));
 sg13g2_tiehi _6811__430 (.L_HI(net614));
 sg13g2_tiehi _6810__431 (.L_HI(net615));
 sg13g2_tiehi _6809__432 (.L_HI(net616));
 sg13g2_tiehi _6808__433 (.L_HI(net617));
 sg13g2_tiehi _6807__434 (.L_HI(net618));
 sg13g2_tiehi _6806__435 (.L_HI(net619));
 sg13g2_tiehi _6805__436 (.L_HI(net620));
 sg13g2_tiehi _6804__437 (.L_HI(net621));
 sg13g2_tiehi _6803__438 (.L_HI(net622));
 sg13g2_tiehi _6802__439 (.L_HI(net623));
 sg13g2_tiehi _6801__440 (.L_HI(net624));
 sg13g2_tiehi _6800__441 (.L_HI(net625));
 sg13g2_tiehi _6799__442 (.L_HI(net626));
 sg13g2_tiehi _6798__443 (.L_HI(net627));
 sg13g2_tiehi _6797__444 (.L_HI(net628));
 sg13g2_tiehi _6796__445 (.L_HI(net629));
 sg13g2_tiehi _6795__446 (.L_HI(net630));
 sg13g2_tiehi _6794__447 (.L_HI(net631));
 sg13g2_tiehi _6793__448 (.L_HI(net632));
 sg13g2_tiehi _6792__449 (.L_HI(net633));
 sg13g2_tiehi _6791__450 (.L_HI(net634));
 sg13g2_tiehi _6790__451 (.L_HI(net635));
 sg13g2_tiehi _6789__452 (.L_HI(net636));
 sg13g2_tiehi _6788__453 (.L_HI(net637));
 sg13g2_tiehi _6787__454 (.L_HI(net638));
 sg13g2_tiehi _6786__455 (.L_HI(net639));
 sg13g2_tiehi _6785__456 (.L_HI(net640));
 sg13g2_tiehi _6784__457 (.L_HI(net641));
 sg13g2_tiehi _6783__458 (.L_HI(net642));
 sg13g2_tiehi _6782__459 (.L_HI(net643));
 sg13g2_tiehi _6781__460 (.L_HI(net644));
 sg13g2_tiehi _6780__461 (.L_HI(net645));
 sg13g2_tiehi _6779__462 (.L_HI(net646));
 sg13g2_tiehi _6778__463 (.L_HI(net647));
 sg13g2_tiehi _6777__464 (.L_HI(net648));
 sg13g2_tiehi _6776__465 (.L_HI(net649));
 sg13g2_tiehi _6775__466 (.L_HI(net650));
 sg13g2_tiehi _6774__467 (.L_HI(net651));
 sg13g2_tiehi _6773__468 (.L_HI(net652));
 sg13g2_tiehi _6772__469 (.L_HI(net653));
 sg13g2_tiehi _6771__470 (.L_HI(net654));
 sg13g2_tiehi _6770__471 (.L_HI(net655));
 sg13g2_tiehi _6769__472 (.L_HI(net656));
 sg13g2_tiehi _6768__473 (.L_HI(net657));
 sg13g2_tiehi _6767__474 (.L_HI(net658));
 sg13g2_tiehi _6766__475 (.L_HI(net659));
 sg13g2_tiehi _6765__476 (.L_HI(net660));
 sg13g2_tiehi _6764__477 (.L_HI(net661));
 sg13g2_tiehi _6763__478 (.L_HI(net662));
 sg13g2_tiehi _6762__479 (.L_HI(net663));
 sg13g2_tiehi _6761__480 (.L_HI(net664));
 sg13g2_tiehi _6760__481 (.L_HI(net665));
 sg13g2_tiehi _6759__482 (.L_HI(net666));
 sg13g2_tiehi _6758__483 (.L_HI(net667));
 sg13g2_tiehi _6757__484 (.L_HI(net668));
 sg13g2_tiehi _6756__485 (.L_HI(net669));
 sg13g2_tiehi _6755__486 (.L_HI(net670));
 sg13g2_tiehi _6754__487 (.L_HI(net671));
 sg13g2_tiehi _6753__488 (.L_HI(net672));
 sg13g2_tiehi _6752__489 (.L_HI(net673));
 sg13g2_tiehi _6751__490 (.L_HI(net674));
 sg13g2_tiehi _6750__491 (.L_HI(net675));
 sg13g2_tiehi _6749__492 (.L_HI(net676));
 sg13g2_tiehi _6748__493 (.L_HI(net677));
 sg13g2_tiehi _6747__494 (.L_HI(net678));
 sg13g2_tiehi _6746__495 (.L_HI(net679));
 sg13g2_tiehi _6745__496 (.L_HI(net680));
 sg13g2_tiehi _6744__497 (.L_HI(net681));
 sg13g2_tiehi _6743__498 (.L_HI(net682));
 sg13g2_tiehi _6742__499 (.L_HI(net683));
 sg13g2_tiehi _6741__500 (.L_HI(net684));
 sg13g2_tiehi _6740__501 (.L_HI(net685));
 sg13g2_tiehi _6739__502 (.L_HI(net686));
 sg13g2_tiehi _6738__503 (.L_HI(net687));
 sg13g2_tiehi _6737__504 (.L_HI(net688));
 sg13g2_tiehi _6736__505 (.L_HI(net689));
 sg13g2_tiehi _6735__506 (.L_HI(net690));
 sg13g2_tiehi _6734__507 (.L_HI(net691));
 sg13g2_tiehi _6733__508 (.L_HI(net692));
 sg13g2_tiehi _6732__509 (.L_HI(net693));
 sg13g2_tiehi _6731__510 (.L_HI(net694));
 sg13g2_tiehi _6730__511 (.L_HI(net695));
 sg13g2_tiehi _6729__512 (.L_HI(net696));
 sg13g2_tiehi _6728__513 (.L_HI(net697));
 sg13g2_tiehi _6727__514 (.L_HI(net698));
 sg13g2_tiehi _6726__515 (.L_HI(net699));
 sg13g2_tiehi _6725__516 (.L_HI(net700));
 sg13g2_tiehi _6724__517 (.L_HI(net701));
 sg13g2_tiehi _6723__518 (.L_HI(net702));
 sg13g2_tiehi _6722__519 (.L_HI(net703));
 sg13g2_tiehi _6721__520 (.L_HI(net704));
 sg13g2_tiehi _6720__521 (.L_HI(net705));
 sg13g2_tiehi _6719__522 (.L_HI(net706));
 sg13g2_tiehi _6718__523 (.L_HI(net707));
 sg13g2_tiehi _6717__524 (.L_HI(net708));
 sg13g2_tiehi _6716__525 (.L_HI(net709));
 sg13g2_tiehi _6715__526 (.L_HI(net710));
 sg13g2_tiehi _6714__527 (.L_HI(net711));
 sg13g2_tiehi _6713__528 (.L_HI(net712));
 sg13g2_tiehi _6712__529 (.L_HI(net713));
 sg13g2_tiehi _6711__530 (.L_HI(net714));
 sg13g2_tiehi _6710__531 (.L_HI(net715));
 sg13g2_tiehi _6709__532 (.L_HI(net716));
 sg13g2_tiehi _6708__533 (.L_HI(net717));
 sg13g2_tiehi _6707__534 (.L_HI(net718));
 sg13g2_tiehi _6706__535 (.L_HI(net719));
 sg13g2_tiehi _6705__536 (.L_HI(net720));
 sg13g2_tiehi _6704__537 (.L_HI(net721));
 sg13g2_tiehi _6703__538 (.L_HI(net722));
 sg13g2_tiehi _6702__539 (.L_HI(net723));
 sg13g2_tiehi _6701__540 (.L_HI(net724));
 sg13g2_tiehi _6391__541 (.L_HI(net725));
 sg13g2_tiehi _6891__542 (.L_HI(net726));
 sg13g2_tiehi _6892__543 (.L_HI(net727));
 sg13g2_tiehi _6893__544 (.L_HI(net728));
 sg13g2_tiehi _6894__545 (.L_HI(net729));
 sg13g2_tiehi _6895__546 (.L_HI(net730));
 sg13g2_tiehi _6896__547 (.L_HI(net731));
 sg13g2_tiehi _6897__548 (.L_HI(net732));
 sg13g2_tiehi _6898__549 (.L_HI(net733));
 sg13g2_tiehi _6899__550 (.L_HI(net734));
 sg13g2_tiehi _6900__551 (.L_HI(net735));
 sg13g2_tiehi _6901__552 (.L_HI(net736));
 sg13g2_tiehi _6902__553 (.L_HI(net737));
 sg13g2_tiehi _6903__554 (.L_HI(net738));
 sg13g2_tiehi _6700__555 (.L_HI(net739));
 sg13g2_tiehi _6699__556 (.L_HI(net740));
 sg13g2_tiehi _6698__557 (.L_HI(net741));
 sg13g2_tiehi _6697__558 (.L_HI(net742));
 sg13g2_tiehi _6696__559 (.L_HI(net743));
 sg13g2_tiehi _6695__560 (.L_HI(net744));
 sg13g2_tiehi _6694__561 (.L_HI(net745));
 sg13g2_tiehi _6693__562 (.L_HI(net746));
 sg13g2_tiehi _6692__563 (.L_HI(net747));
 sg13g2_tiehi _6691__564 (.L_HI(net748));
 sg13g2_tiehi _6690__565 (.L_HI(net749));
 sg13g2_tiehi _6689__566 (.L_HI(net750));
 sg13g2_tiehi _6688__567 (.L_HI(net751));
 sg13g2_tiehi _6687__568 (.L_HI(net752));
 sg13g2_tiehi _6686__569 (.L_HI(net753));
 sg13g2_tiehi _6685__570 (.L_HI(net754));
 sg13g2_tiehi _6684__571 (.L_HI(net755));
 sg13g2_tiehi _6683__572 (.L_HI(net756));
 sg13g2_tiehi heichips25_CORDIC_573 (.L_HI(net757));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo heichips25_CORDIC_25 (.L_LO(net25));
 sg13g2_tielo heichips25_CORDIC_26 (.L_LO(net26));
 sg13g2_tielo heichips25_CORDIC_27 (.L_LO(net27));
 sg13g2_tielo heichips25_CORDIC_28 (.L_LO(net28));
 sg13g2_tielo heichips25_CORDIC_29 (.L_LO(net29));
 sg13g2_tielo heichips25_CORDIC_30 (.L_LO(net30));
 sg13g2_tielo heichips25_CORDIC_31 (.L_LO(net31));
 sg13g2_tielo heichips25_CORDIC_32 (.L_LO(net32));
 sg13g2_tielo heichips25_CORDIC_33 (.L_LO(net33));
 sg13g2_tielo heichips25_CORDIC_34 (.L_LO(net34));
 sg13g2_tielo heichips25_CORDIC_35 (.L_LO(net35));
 sg13g2_tielo heichips25_CORDIC_36 (.L_LO(net36));
 sg13g2_tielo heichips25_CORDIC_37 (.L_LO(net37));
 sg13g2_tielo heichips25_CORDIC_38 (.L_LO(net38));
 sg13g2_tielo heichips25_CORDIC_39 (.L_LO(net39));
 sg13g2_tiehi _6682__40 (.L_HI(net40));
 sg13g2_buf_1 _7474_ (.A(pwm_data),
    .X(net17));
 sg13g2_buf_1 _7475_ (.A(net21),
    .X(net18));
 sg13g2_buf_1 _7476_ (.A(net22),
    .X(net19));
 sg13g2_buf_1 _7477_ (.A(\u_angle_cordic_12b_pmod.u_vga_top.vsync ),
    .X(net20));
 sg13g2_buf_1 _7478_ (.A(hsync_sig),
    .X(net23));
 sg13g2_buf_8 fanout372 (.A(net373),
    .X(net372));
 sg13g2_buf_8 fanout373 (.A(_0991_),
    .X(net373));
 sg13g2_buf_8 fanout374 (.A(net375),
    .X(net374));
 sg13g2_buf_8 fanout375 (.A(_0989_),
    .X(net375));
 sg13g2_buf_8 fanout376 (.A(net377),
    .X(net376));
 sg13g2_buf_8 fanout377 (.A(net378),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_0988_),
    .X(net378));
 sg13g2_buf_8 fanout379 (.A(_2007_),
    .X(net379));
 sg13g2_buf_8 fanout380 (.A(_1934_),
    .X(net380));
 sg13g2_buf_8 fanout381 (.A(_1233_),
    .X(net381));
 sg13g2_buf_8 fanout382 (.A(net383),
    .X(net382));
 sg13g2_buf_8 fanout383 (.A(_1159_),
    .X(net383));
 sg13g2_buf_8 fanout384 (.A(net385),
    .X(net384));
 sg13g2_buf_8 fanout385 (.A(_1416_),
    .X(net385));
 sg13g2_buf_8 fanout386 (.A(net387),
    .X(net386));
 sg13g2_buf_8 fanout387 (.A(_1342_),
    .X(net387));
 sg13g2_buf_8 fanout388 (.A(net390),
    .X(net388));
 sg13g2_buf_8 fanout389 (.A(net390),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_1722_),
    .X(net390));
 sg13g2_buf_8 fanout391 (.A(net392),
    .X(net391));
 sg13g2_buf_8 fanout392 (.A(_1660_),
    .X(net392));
 sg13g2_buf_8 fanout393 (.A(net394),
    .X(net393));
 sg13g2_buf_8 fanout394 (.A(_1522_),
    .X(net394));
 sg13g2_buf_8 fanout395 (.A(_1843_),
    .X(net395));
 sg13g2_buf_8 fanout396 (.A(_1842_),
    .X(net396));
 sg13g2_buf_8 fanout397 (.A(net398),
    .X(net397));
 sg13g2_buf_8 fanout398 (.A(net399),
    .X(net398));
 sg13g2_buf_8 fanout399 (.A(_1783_),
    .X(net399));
 sg13g2_buf_8 fanout400 (.A(net401),
    .X(net400));
 sg13g2_buf_8 fanout401 (.A(_1592_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_2857_),
    .X(net402));
 sg13g2_buf_8 fanout403 (.A(_0647_),
    .X(net403));
 sg13g2_buf_8 fanout404 (.A(_0646_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_0646_),
    .X(net405));
 sg13g2_buf_8 fanout406 (.A(_0644_),
    .X(net406));
 sg13g2_buf_8 fanout407 (.A(_0643_),
    .X(net407));
 sg13g2_buf_8 fanout408 (.A(_0642_),
    .X(net408));
 sg13g2_buf_8 fanout409 (.A(_0641_),
    .X(net409));
 sg13g2_buf_8 fanout410 (.A(net411),
    .X(net410));
 sg13g2_buf_8 fanout411 (.A(_0600_),
    .X(net411));
 sg13g2_buf_8 fanout412 (.A(_0592_),
    .X(net412));
 sg13g2_buf_8 fanout413 (.A(_0573_),
    .X(net413));
 sg13g2_buf_1 fanout414 (.A(_0573_),
    .X(net414));
 sg13g2_buf_8 fanout415 (.A(_0564_),
    .X(net415));
 sg13g2_buf_8 fanout416 (.A(_0562_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_0562_),
    .X(net417));
 sg13g2_buf_8 fanout418 (.A(_0553_),
    .X(net418));
 sg13g2_buf_8 fanout419 (.A(net423),
    .X(net419));
 sg13g2_buf_8 fanout420 (.A(net423),
    .X(net420));
 sg13g2_buf_8 fanout421 (.A(net422),
    .X(net421));
 sg13g2_buf_8 fanout422 (.A(net423),
    .X(net422));
 sg13g2_buf_8 fanout423 (.A(net440),
    .X(net423));
 sg13g2_buf_8 fanout424 (.A(net428),
    .X(net424));
 sg13g2_buf_8 fanout425 (.A(net428),
    .X(net425));
 sg13g2_buf_8 fanout426 (.A(net428),
    .X(net426));
 sg13g2_buf_1 fanout427 (.A(net428),
    .X(net427));
 sg13g2_buf_8 fanout428 (.A(net440),
    .X(net428));
 sg13g2_buf_8 fanout429 (.A(net434),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(net434),
    .X(net430));
 sg13g2_buf_8 fanout431 (.A(net434),
    .X(net431));
 sg13g2_buf_8 fanout432 (.A(net434),
    .X(net432));
 sg13g2_buf_8 fanout433 (.A(net434),
    .X(net433));
 sg13g2_buf_8 fanout434 (.A(net440),
    .X(net434));
 sg13g2_buf_8 fanout435 (.A(net438),
    .X(net435));
 sg13g2_buf_8 fanout436 (.A(net437),
    .X(net436));
 sg13g2_buf_8 fanout437 (.A(net438),
    .X(net437));
 sg13g2_buf_8 fanout438 (.A(net439),
    .X(net438));
 sg13g2_buf_8 fanout439 (.A(net440),
    .X(net439));
 sg13g2_buf_8 fanout440 (.A(_0546_),
    .X(net440));
 sg13g2_buf_8 fanout441 (.A(net443),
    .X(net441));
 sg13g2_buf_1 fanout442 (.A(net443),
    .X(net442));
 sg13g2_buf_8 fanout443 (.A(net451),
    .X(net443));
 sg13g2_buf_8 fanout444 (.A(net447),
    .X(net444));
 sg13g2_buf_8 fanout445 (.A(net447),
    .X(net445));
 sg13g2_buf_1 fanout446 (.A(net447),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(net451),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(net449),
    .X(net448));
 sg13g2_buf_8 fanout449 (.A(net450),
    .X(net449));
 sg13g2_buf_8 fanout450 (.A(net451),
    .X(net450));
 sg13g2_buf_8 fanout451 (.A(net851),
    .X(net451));
 sg13g2_buf_8 fanout452 (.A(net456),
    .X(net452));
 sg13g2_buf_1 fanout453 (.A(net456),
    .X(net453));
 sg13g2_buf_8 fanout454 (.A(net456),
    .X(net454));
 sg13g2_buf_1 fanout455 (.A(net456),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(net473),
    .X(net456));
 sg13g2_buf_8 fanout457 (.A(net458),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(net461),
    .X(net458));
 sg13g2_buf_8 fanout459 (.A(net461),
    .X(net459));
 sg13g2_buf_1 fanout460 (.A(net461),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(net473),
    .X(net461));
 sg13g2_buf_8 fanout462 (.A(net466),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(net465),
    .X(net463));
 sg13g2_buf_8 fanout464 (.A(net465),
    .X(net464));
 sg13g2_buf_8 fanout465 (.A(net466),
    .X(net465));
 sg13g2_buf_8 fanout466 (.A(net473),
    .X(net466));
 sg13g2_buf_8 fanout467 (.A(net468),
    .X(net467));
 sg13g2_buf_8 fanout468 (.A(net472),
    .X(net468));
 sg13g2_buf_8 fanout469 (.A(net471),
    .X(net469));
 sg13g2_buf_1 fanout470 (.A(net471),
    .X(net470));
 sg13g2_buf_8 fanout471 (.A(net472),
    .X(net471));
 sg13g2_buf_8 fanout472 (.A(net473),
    .X(net472));
 sg13g2_buf_8 fanout473 (.A(net851),
    .X(net473));
 sg13g2_buf_8 fanout474 (.A(net476),
    .X(net474));
 sg13g2_buf_1 fanout475 (.A(net476),
    .X(net475));
 sg13g2_buf_8 fanout476 (.A(net491),
    .X(net476));
 sg13g2_buf_8 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_8 fanout478 (.A(net480),
    .X(net478));
 sg13g2_buf_8 fanout479 (.A(net480),
    .X(net479));
 sg13g2_buf_8 fanout480 (.A(net491),
    .X(net480));
 sg13g2_buf_8 fanout481 (.A(net482),
    .X(net481));
 sg13g2_buf_1 fanout482 (.A(net490),
    .X(net482));
 sg13g2_buf_8 fanout483 (.A(net485),
    .X(net483));
 sg13g2_buf_1 fanout484 (.A(net485),
    .X(net484));
 sg13g2_buf_8 fanout485 (.A(net490),
    .X(net485));
 sg13g2_buf_8 fanout486 (.A(net487),
    .X(net486));
 sg13g2_buf_1 fanout487 (.A(net490),
    .X(net487));
 sg13g2_buf_8 fanout488 (.A(net490),
    .X(net488));
 sg13g2_buf_1 fanout489 (.A(net490),
    .X(net489));
 sg13g2_buf_8 fanout490 (.A(net491),
    .X(net490));
 sg13g2_buf_8 fanout491 (.A(net505),
    .X(net491));
 sg13g2_buf_8 fanout492 (.A(net494),
    .X(net492));
 sg13g2_buf_1 fanout493 (.A(net494),
    .X(net493));
 sg13g2_buf_1 fanout494 (.A(net495),
    .X(net494));
 sg13g2_buf_1 fanout495 (.A(net505),
    .X(net495));
 sg13g2_buf_8 fanout496 (.A(net500),
    .X(net496));
 sg13g2_buf_1 fanout497 (.A(net500),
    .X(net497));
 sg13g2_buf_8 fanout498 (.A(net500),
    .X(net498));
 sg13g2_buf_1 fanout499 (.A(net500),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(net505),
    .X(net500));
 sg13g2_buf_8 fanout501 (.A(net504),
    .X(net501));
 sg13g2_buf_8 fanout502 (.A(net504),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(net504),
    .X(net503));
 sg13g2_buf_8 fanout504 (.A(net505),
    .X(net504));
 sg13g2_buf_8 fanout505 (.A(net851),
    .X(net505));
 sg13g2_buf_8 fanout506 (.A(net939),
    .X(net506));
 sg13g2_buf_8 fanout507 (.A(net511),
    .X(net507));
 sg13g2_buf_8 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(net511),
    .X(net509));
 sg13g2_buf_8 fanout510 (.A(net511),
    .X(net510));
 sg13g2_buf_8 fanout511 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].z_sign ),
    .X(net511));
 sg13g2_buf_8 fanout512 (.A(net514),
    .X(net512));
 sg13g2_buf_8 fanout513 (.A(net514),
    .X(net513));
 sg13g2_buf_8 fanout514 (.A(net1247),
    .X(net514));
 sg13g2_buf_8 fanout515 (.A(net516),
    .X(net515));
 sg13g2_buf_8 fanout516 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].z_sign ),
    .X(net516));
 sg13g2_buf_8 fanout517 (.A(net518),
    .X(net517));
 sg13g2_buf_8 fanout518 (.A(net519),
    .X(net518));
 sg13g2_buf_8 fanout519 (.A(net520),
    .X(net519));
 sg13g2_buf_8 fanout520 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].z_sign ),
    .X(net520));
 sg13g2_buf_8 fanout521 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].z_sign ),
    .X(net521));
 sg13g2_buf_1 fanout522 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].z_sign ),
    .X(net522));
 sg13g2_buf_8 fanout523 (.A(net525),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(net525),
    .X(net524));
 sg13g2_buf_8 fanout525 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].z_sign ),
    .X(net525));
 sg13g2_buf_8 fanout526 (.A(net530),
    .X(net526));
 sg13g2_buf_1 fanout527 (.A(net530),
    .X(net527));
 sg13g2_buf_8 fanout528 (.A(net530),
    .X(net528));
 sg13g2_buf_1 fanout529 (.A(net530),
    .X(net529));
 sg13g2_buf_8 fanout530 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].z_sign ),
    .X(net530));
 sg13g2_buf_8 fanout531 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].z_sign ),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].z_sign ),
    .X(net532));
 sg13g2_buf_8 fanout533 (.A(net534),
    .X(net533));
 sg13g2_buf_8 fanout534 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].z_sign ),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.sqr_amp[0] ),
    .X(net535));
 sg13g2_buf_8 fanout536 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].z_sign ),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(net538),
    .X(net537));
 sg13g2_buf_1 fanout538 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].z_sign ),
    .X(net538));
 sg13g2_buf_8 fanout539 (.A(net540),
    .X(net539));
 sg13g2_buf_8 fanout540 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].z_sign ),
    .X(net540));
 sg13g2_buf_8 fanout541 (.A(net542),
    .X(net541));
 sg13g2_buf_8 fanout542 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].z_sign ),
    .X(net542));
 sg13g2_buf_8 fanout543 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].z_sign ),
    .X(net543));
 sg13g2_buf_8 fanout544 (.A(net545),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(\u_angle_cordic_12b_pmod.waveform_sel_reg[1] ),
    .X(net545));
 sg13g2_buf_8 fanout546 (.A(net547),
    .X(net546));
 sg13g2_buf_8 fanout547 (.A(\u_angle_cordic_12b_pmod.waveform_sel_reg[0] ),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(net551),
    .X(net548));
 sg13g2_buf_8 fanout549 (.A(net551),
    .X(net549));
 sg13g2_buf_1 fanout550 (.A(net551),
    .X(net550));
 sg13g2_buf_1 fanout551 (.A(net1179),
    .X(net551));
 sg13g2_buf_8 fanout552 (.A(\u_angle_cordic_12b_pmod.u_vga_top.pixel_clk_en ),
    .X(net552));
 sg13g2_buf_8 fanout553 (.A(net554),
    .X(net553));
 sg13g2_buf_8 fanout554 (.A(\u_angle_cordic_12b_pmod.u_vga_top.pixel_clk_en ),
    .X(net554));
 sg13g2_buf_8 fanout555 (.A(net1043),
    .X(net555));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[1]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[2]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[3]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[4]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[5]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[6]),
    .X(net16));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[7]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[0]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[1]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[3]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[4]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[5]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[7]));
 sg13g2_tielo heichips25_CORDIC_24 (.L_LO(net24));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_4_5_0_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_4_6_0_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_4_7_0_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_4_9_0_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_4_10_0_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_4_11_0_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_4_12_0_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_4_13_0_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_4_14_0_clk));
 sg13g2_buf_8 clkload12 (.A(clknet_4_15_0_clk));
 sg13g2_buf_8 clkload13 (.A(clknet_leaf_66_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][9] ),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold2 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][1] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold3 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][0] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold4 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][0] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0440_),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold6 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[0] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold7 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][2] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold8 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][0] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold9 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][2] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold10 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][1] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold11 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][1] ),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold12 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][3] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold13 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][0] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold14 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][6] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold15 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][0] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold16 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][4] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold17 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][1] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold18 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][5] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold19 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][7] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0050_),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold21 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][7] ),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold22 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][2] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold23 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][8] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold24 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][6] ),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0049_),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold26 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][3] ),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold27 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][3] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold28 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][8] ),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold29 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][4] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold30 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][6] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold31 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][9] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold32 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][10] ),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold33 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][2] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold34 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][0] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold35 (.A(\u_angle_cordic_12b_pmod.u_vga_top.clk_div_cnt[0] ),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold36 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][4] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold37 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][9] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold38 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][10] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold39 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][7] ),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0496_),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold41 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][0] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold42 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][1] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold43 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][0] ),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold44 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][5] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold45 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][1] ),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold46 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[11] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold47 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][2] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold48 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][4] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold49 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][0] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold50 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][8] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold51 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][5] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold52 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][0] ),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold53 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][5] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold54 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][10] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0337_),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold56 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[10] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0006_),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold58 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[0][10] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0488_),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold60 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][1] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold61 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][10] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold62 (.A(_0132_),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold63 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][3] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold64 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[8] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold65 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.x_start[0] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0003_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold67 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[5] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold68 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[11][11] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold69 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][10] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0375_),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold71 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[7] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0077_),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold73 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][1] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold74 (.A(\u_angle_cordic_12b_pmod.u_vga_top.clk_div_cnt[1] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold75 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][10] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0170_),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold77 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][2] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold78 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[9] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0005_),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold80 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][10] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0299_),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold82 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[11][11] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold83 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[1] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold84 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][6] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold85 (.A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[8] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0028_),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold87 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[5] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0506_),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold89 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[4] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold90 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[9] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0510_),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold92 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[3] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0524_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold94 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.resetn ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold95 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][0] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0327_),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold97 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[15] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0516_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold99 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[6] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold100 (.A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[0] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0020_),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold102 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[10] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0635_),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0002_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold105 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][3] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold106 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[10] ),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0041_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold108 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[9] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold109 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[6] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0857_),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0017_),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold112 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[7] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0868_),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0018_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold115 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[10] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0183_),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold117 (.A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[1] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0875_),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0021_),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold120 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][1] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold121 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[11] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold122 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[0] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold123 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[10] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold124 (.A(_2914_),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold125 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[0] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0848_),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0012_),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold128 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[7] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0063_),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold130 (.A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[9] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0893_),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold132 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[8] ),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0872_),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0019_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold135 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[2] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0852_),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0014_),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold138 (.A(net21),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0820_),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0009_),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold141 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[2] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold142 (.A(_2900_),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0503_),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold144 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[7] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0038_),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold146 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[10] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold147 (.A(_2428_),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0363_),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold149 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[1] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0849_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0013_),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold152 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[3] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0853_),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0015_),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold155 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][0] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold156 (.A(_1962_),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold157 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[8] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0920_),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold159 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[16] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold160 (.A(_2924_),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold161 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[8] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold162 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle[2] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold163 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[2] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0033_),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold165 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][0] ),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold166 (.A(_1305_),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold167 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[1] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0057_),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold169 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[4] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold170 (.A(_2904_),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0505_),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold172 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[5] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0004_),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold174 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[3] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold175 (.A(_2902_),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold176 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][0] ),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold177 (.A(_2269_),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0338_),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold179 (.A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[3] ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0879_),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0023_),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold182 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[0].z_sign ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold183 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[0] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold184 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[6] ),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0917_),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0037_),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold187 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_pos[4] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0016_),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold189 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][0] ),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold190 (.A(_1770_),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold191 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[4] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0060_),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold193 (.A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[2] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0877_),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold195 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[6] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0062_),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold197 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[3] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0059_),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold199 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[8] ),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold200 (.A(_2911_),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold201 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[13] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold202 (.A(_2920_),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0514_),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold204 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[5] ),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold205 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][0] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold206 (.A(_1188_),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0108_),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold208 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][1] ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold209 (.A(_2736_),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold210 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[0].y_shr[0] ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold211 (.A(_2858_),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0452_),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold213 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][0] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold214 (.A(_2072_),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0300_),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold216 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[2][0] ),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold217 (.A(_2555_),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold218 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[11] ),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold219 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][0] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold220 (.A(_1492_),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold221 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[3] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0034_),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold223 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[2] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold224 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[12] ),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold225 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[10] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold226 (.A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[10] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0030_),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold228 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][0] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold229 (.A(_1378_),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0146_),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold231 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][0] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold232 (.A(_1826_),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0236_),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold234 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[0] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0109_),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold236 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][0] ),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold237 (.A(_1563_),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0184_),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold239 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[0] ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0147_),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold241 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][0] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold242 (.A(_1703_),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0211_),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold244 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[9] ),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0040_),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold246 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[4] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0913_),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold248 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][2] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold249 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][1] ),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold250 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[1] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold251 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[0] ),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0301_),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold253 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[3][0] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold254 (.A(_2350_),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold255 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.tri_amp[9] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0065_),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold257 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][0] ),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold258 (.A(_2474_),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold259 (.A(_0376_),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold260 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[0] ),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0185_),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold262 (.A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[7] ),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0891_),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0027_),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold265 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[14] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold266 (.A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[4] ),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold267 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[1] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0032_),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold269 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][2] ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold270 (.A(_1265_),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0123_),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold272 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[17] ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold273 (.A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[6] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0889_),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0026_),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold276 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][0] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold277 (.A(_1884_),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0262_),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold279 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][10] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold280 (.A(_1114_),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold281 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][4] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0163_),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold283 (.A(\u_angle_cordic_12b_pmod.u_vga_top.h_cnt[5] ),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold284 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[0][0] ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0469_),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold286 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[0].y_shr[10] ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold287 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[0] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold288 (.A(_0212_),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold289 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][0] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold290 (.A(_2653_),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0414_),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold292 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][3] ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0444_),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold294 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][7] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold295 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[0] ),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0237_),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold297 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[4][0] ),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold298 (.A(_2150_),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold299 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[5] ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold300 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][3] ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold301 (.A(_1079_),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0086_),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold303 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][5] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0088_),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold305 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][1] ),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold306 (.A(_1966_),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0276_),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold308 (.A(net22),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0830_),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0010_),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold311 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][10] ),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold312 (.A(_2651_),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold313 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[0].y_shr[11] ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold314 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][8] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold315 (.A(_2848_),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0449_),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold317 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][2] ),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0328_),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold319 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[0] ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold320 (.A(_0415_),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold321 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][7] ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0371_),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold323 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][4] ),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0125_),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold325 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][0] ),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold326 (.A(_1638_),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold327 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][5] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0369_),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold329 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][8] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold330 (.A(_1481_),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold331 (.A(_0167_),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold332 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][3] ),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0330_),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold334 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][6] ),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0205_),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold336 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[0] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0903_),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold338 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][4] ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0292_),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold340 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][1] ),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0134_),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold342 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][10] ),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold343 (.A(_2856_),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold344 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[0] ),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0263_),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold346 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][0] ),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold347 (.A(_1115_),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0096_),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold349 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][6] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold350 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[7] ),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold351 (.A(_2909_),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0508_),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold353 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][8] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0129_),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold355 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][4] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0229_),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold357 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.cnt[6] ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold358 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][9] ),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0092_),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold360 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[8] ),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold361 (.A(_2423_),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0362_),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold363 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][5] ),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold364 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][9] ),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold365 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][6] ),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0231_),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold367 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][8] ),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold368 (.A(_2265_),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold369 (.A(_0336_),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold370 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][9] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold371 (.A(_2470_),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0374_),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold373 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][11] ),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold374 (.A(_2726_),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold375 (.A(_0426_),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold376 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][7] ),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold377 (.A(_1474_),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold378 (.A(_1476_),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold379 (.A(_0166_),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold380 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][8] ),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold381 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][7] ),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold382 (.A(_1287_),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold383 (.A(_1289_),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold384 (.A(_0128_),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold385 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[9][10] ),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0197_),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold387 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][6] ),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0294_),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold389 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[2][1] ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold390 (.A(_2559_),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0390_),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold392 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][8] ),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold393 (.A(_1101_),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold394 (.A(_1103_),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold395 (.A(_0091_),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold396 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][5] ),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold397 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][9] ),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold398 (.A(_0411_),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold399 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][7] ),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold400 (.A(_0333_),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold401 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[3] ),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold402 (.A(_0144_),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold403 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][1] ),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0225_),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold405 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][6] ),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold406 (.A(_1926_),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold407 (.A(_0268_),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold408 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][1] ),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0172_),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold410 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][4] ),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold411 (.A(_0216_),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold412 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][10] ),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0157_),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold414 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][9] ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold415 (.A(_2263_),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold416 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][8] ),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0220_),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold418 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][7] ),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0090_),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold420 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[3] ),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0182_),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold422 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.angle_gen.up ),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0055_),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold424 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[3] ),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold425 (.A(_0284_),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold426 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[2] ),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0104_),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold428 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][9] ),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold429 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][9] ),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0233_),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold431 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[1] ),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold432 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][7] ),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold433 (.A(_1537_),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold434 (.A(_0178_),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold435 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][6] ),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold436 (.A(_0127_),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold437 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][11] ),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold438 (.A(_0349_),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold439 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[10].y_shr[1] ),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold440 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][11] ),
    .X(net1197));
 sg13g2_dlygate4sd3_1 hold441 (.A(_0247_),
    .X(net1198));
 sg13g2_dlygate4sd3_1 hold442 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][12] ),
    .X(net1199));
 sg13g2_dlygate4sd3_1 hold443 (.A(_0120_),
    .X(net1200));
 sg13g2_dlygate4sd3_1 hold444 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[2] ),
    .X(net1201));
 sg13g2_dlygate4sd3_1 hold445 (.A(_1698_),
    .X(net1202));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0210_),
    .X(net1203));
 sg13g2_dlygate4sd3_1 hold447 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][4] ),
    .X(net1204));
 sg13g2_dlygate4sd3_1 hold448 (.A(_0368_),
    .X(net1205));
 sg13g2_dlygate4sd3_1 hold449 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][3] ),
    .X(net1206));
 sg13g2_dlygate4sd3_1 hold450 (.A(_0149_),
    .X(net1207));
 sg13g2_dlygate4sd3_1 hold451 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[1] ),
    .X(net1208));
 sg13g2_dlygate4sd3_1 hold452 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][5] ),
    .X(net1209));
 sg13g2_dlygate4sd3_1 hold453 (.A(_2687_),
    .X(net1210));
 sg13g2_dlygate4sd3_1 hold454 (.A(_0419_),
    .X(net1211));
 sg13g2_dlygate4sd3_1 hold455 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][4] ),
    .X(net1212));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0175_),
    .X(net1213));
 sg13g2_dlygate4sd3_1 hold457 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][6] ),
    .X(net1214));
 sg13g2_dlygate4sd3_1 hold458 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][12] ),
    .X(net1215));
 sg13g2_dlygate4sd3_1 hold459 (.A(_0223_),
    .X(net1216));
 sg13g2_dlygate4sd3_1 hold460 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][12] ),
    .X(net1217));
 sg13g2_dlygate4sd3_1 hold461 (.A(_0388_),
    .X(net1218));
 sg13g2_dlygate4sd3_1 hold462 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][8] ),
    .X(net1219));
 sg13g2_dlygate4sd3_1 hold463 (.A(_1870_),
    .X(net1220));
 sg13g2_dlygate4sd3_1 hold464 (.A(_0244_),
    .X(net1221));
 sg13g2_dlygate4sd3_1 hold465 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][6] ),
    .X(net1222));
 sg13g2_dlygate4sd3_1 hold466 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][2] ),
    .X(net1223));
 sg13g2_dlygate4sd3_1 hold467 (.A(_1390_),
    .X(net1224));
 sg13g2_dlygate4sd3_1 hold468 (.A(_1391_),
    .X(net1225));
 sg13g2_dlygate4sd3_1 hold469 (.A(_0148_),
    .X(net1226));
 sg13g2_dlygate4sd3_1 hold470 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[5] ),
    .X(net1227));
 sg13g2_dlygate4sd3_1 hold471 (.A(_2030_),
    .X(net1228));
 sg13g2_dlygate4sd3_1 hold472 (.A(_0286_),
    .X(net1229));
 sg13g2_dlygate4sd3_1 hold473 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[0] ),
    .X(net1230));
 sg13g2_dlygate4sd3_1 hold474 (.A(_2275_),
    .X(net1231));
 sg13g2_dlygate4sd3_1 hold475 (.A(_0339_),
    .X(net1232));
 sg13g2_dlygate4sd3_1 hold476 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][12] ),
    .X(net1233));
 sg13g2_dlygate4sd3_1 hold477 (.A(_0312_),
    .X(net1234));
 sg13g2_dlygate4sd3_1 hold478 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][6] ),
    .X(net1235));
 sg13g2_dlygate4sd3_1 hold479 (.A(_0446_),
    .X(net1236));
 sg13g2_dlygate4sd3_1 hold480 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][4] ),
    .X(net1237));
 sg13g2_dlygate4sd3_1 hold481 (.A(_1666_),
    .X(net1238));
 sg13g2_dlygate4sd3_1 hold482 (.A(_0203_),
    .X(net1239));
 sg13g2_dlygate4sd3_1 hold483 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[3][1] ),
    .X(net1240));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0352_),
    .X(net1241));
 sg13g2_dlygate4sd3_1 hold485 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[0] ),
    .X(net1242));
 sg13g2_dlygate4sd3_1 hold486 (.A(_2480_),
    .X(net1243));
 sg13g2_dlygate4sd3_1 hold487 (.A(_0377_),
    .X(net1244));
 sg13g2_dlygate4sd3_1 hold488 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][3] ),
    .X(net1245));
 sg13g2_dlygate4sd3_1 hold489 (.A(_0278_),
    .X(net1246));
 sg13g2_dlygate4sd3_1 hold490 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].z_sign ),
    .X(net1247));
 sg13g2_dlygate4sd3_1 hold491 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[2] ),
    .X(net1248));
 sg13g2_dlygate4sd3_1 hold492 (.A(_2580_),
    .X(net1249));
 sg13g2_dlygate4sd3_1 hold493 (.A(_0393_),
    .X(net1250));
 sg13g2_dlygate4sd3_1 hold494 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][6] ),
    .X(net1251));
 sg13g2_dlygate4sd3_1 hold495 (.A(_0218_),
    .X(net1252));
 sg13g2_dlygate4sd3_1 hold496 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][6] ),
    .X(net1253));
 sg13g2_dlygate4sd3_1 hold497 (.A(_0177_),
    .X(net1254));
 sg13g2_dlygate4sd3_1 hold498 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][3] ),
    .X(net1255));
 sg13g2_dlygate4sd3_1 hold499 (.A(_2090_),
    .X(net1256));
 sg13g2_dlygate4sd3_1 hold500 (.A(_0303_),
    .X(net1257));
 sg13g2_dlygate4sd3_1 hold501 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][12] ),
    .X(net1258));
 sg13g2_dlygate4sd3_1 hold502 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][7] ),
    .X(net1259));
 sg13g2_dlygate4sd3_1 hold503 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][9] ),
    .X(net1260));
 sg13g2_dlygate4sd3_1 hold504 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[1] ),
    .X(net1261));
 sg13g2_dlygate4sd3_1 hold505 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][12] ),
    .X(net1262));
 sg13g2_dlygate4sd3_1 hold506 (.A(_0158_),
    .X(net1263));
 sg13g2_dlygate4sd3_1 hold507 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][2] ),
    .X(net1264));
 sg13g2_dlygate4sd3_1 hold508 (.A(_2738_),
    .X(net1265));
 sg13g2_dlygate4sd3_1 hold509 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[6][4] ),
    .X(net1266));
 sg13g2_dlygate4sd3_1 hold510 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][7] ),
    .X(net1267));
 sg13g2_dlygate4sd3_1 hold511 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][9] ),
    .X(net1268));
 sg13g2_dlygate4sd3_1 hold512 (.A(_2065_),
    .X(net1269));
 sg13g2_dlygate4sd3_1 hold513 (.A(_0297_),
    .X(net1270));
 sg13g2_dlygate4sd3_1 hold514 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][5] ),
    .X(net1271));
 sg13g2_dlygate4sd3_1 hold515 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][2] ),
    .X(net1272));
 sg13g2_dlygate4sd3_1 hold516 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][10] ),
    .X(net1273));
 sg13g2_dlygate4sd3_1 hold517 (.A(_0195_),
    .X(net1274));
 sg13g2_dlygate4sd3_1 hold518 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][4] ),
    .X(net1275));
 sg13g2_dlygate4sd3_1 hold519 (.A(_0267_),
    .X(net1276));
 sg13g2_dlygate4sd3_1 hold520 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][2] ),
    .X(net1277));
 sg13g2_dlygate4sd3_1 hold521 (.A(_1198_),
    .X(net1278));
 sg13g2_dlygate4sd3_1 hold522 (.A(_1199_),
    .X(net1279));
 sg13g2_dlygate4sd3_1 hold523 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][2] ),
    .X(net1280));
 sg13g2_dlygate4sd3_1 hold524 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[11] ),
    .X(net1281));
 sg13g2_dlygate4sd3_1 hold525 (.A(_2817_),
    .X(net1282));
 sg13g2_dlygate4sd3_1 hold526 (.A(_0439_),
    .X(net1283));
 sg13g2_dlygate4sd3_1 hold527 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[7][3] ),
    .X(net1284));
 sg13g2_dlygate4sd3_1 hold528 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[10] ),
    .X(net1285));
 sg13g2_dlygate4sd3_1 hold529 (.A(_0325_),
    .X(net1286));
 sg13g2_dlygate4sd3_1 hold530 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[10] ),
    .X(net1287));
 sg13g2_dlygate4sd3_1 hold531 (.A(_0145_),
    .X(net1288));
 sg13g2_dlygate4sd3_1 hold532 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][9] ),
    .X(net1289));
 sg13g2_dlygate4sd3_1 hold533 (.A(_0271_),
    .X(net1290));
 sg13g2_dlygate4sd3_1 hold534 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][11] ),
    .X(net1291));
 sg13g2_dlygate4sd3_1 hold535 (.A(_0273_),
    .X(net1292));
 sg13g2_dlygate4sd3_1 hold536 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][5] ),
    .X(net1293));
 sg13g2_dlygate4sd3_1 hold537 (.A(_0189_),
    .X(net1294));
 sg13g2_dlygate4sd3_1 hold538 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][4] ),
    .X(net1295));
 sg13g2_dlygate4sd3_1 hold539 (.A(_2680_),
    .X(net1296));
 sg13g2_dlygate4sd3_1 hold540 (.A(_0418_),
    .X(net1297));
 sg13g2_dlygate4sd3_1 hold541 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[2] ),
    .X(net1298));
 sg13g2_dlygate4sd3_1 hold542 (.A(_0430_),
    .X(net1299));
 sg13g2_dlygate4sd3_1 hold543 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[4] ),
    .X(net1300));
 sg13g2_dlygate4sd3_1 hold544 (.A(_0106_),
    .X(net1301));
 sg13g2_dlygate4sd3_1 hold545 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][2] ),
    .X(net1302));
 sg13g2_dlygate4sd3_1 hold546 (.A(_0340_),
    .X(net1303));
 sg13g2_dlygate4sd3_1 hold547 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[4][1] ),
    .X(net1304));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0314_),
    .X(net1305));
 sg13g2_dlygate4sd3_1 hold549 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][6] ),
    .X(net1306));
 sg13g2_dlygate4sd3_1 hold550 (.A(_2516_),
    .X(net1307));
 sg13g2_dlygate4sd3_1 hold551 (.A(_0382_),
    .X(net1308));
 sg13g2_dlygate4sd3_1 hold552 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[10] ),
    .X(net1309));
 sg13g2_dlygate4sd3_1 hold553 (.A(_0107_),
    .X(net1310));
 sg13g2_dlygate4sd3_1 hold554 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][3] ),
    .X(net1311));
 sg13g2_dlygate4sd3_1 hold555 (.A(_0187_),
    .X(net1312));
 sg13g2_dlygate4sd3_1 hold556 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][8] ),
    .X(net1313));
 sg13g2_dlygate4sd3_1 hold557 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[6] ),
    .X(net1314));
 sg13g2_dlygate4sd3_1 hold558 (.A(_2033_),
    .X(net1315));
 sg13g2_dlygate4sd3_1 hold559 (.A(_0287_),
    .X(net1316));
 sg13g2_dlygate4sd3_1 hold560 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[1] ),
    .X(net1317));
 sg13g2_dlygate4sd3_1 hold561 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][7] ),
    .X(net1318));
 sg13g2_dlygate4sd3_1 hold562 (.A(_2700_),
    .X(net1319));
 sg13g2_dlygate4sd3_1 hold563 (.A(_2710_),
    .X(net1320));
 sg13g2_dlygate4sd3_1 hold564 (.A(_0422_),
    .X(net1321));
 sg13g2_dlygate4sd3_1 hold565 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][3] ),
    .X(net1322));
 sg13g2_dlygate4sd3_1 hold566 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[10] ),
    .X(net1323));
 sg13g2_dlygate4sd3_1 hold567 (.A(_0401_),
    .X(net1324));
 sg13g2_dlygate4sd3_1 hold568 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[2][8] ),
    .X(net1325));
 sg13g2_dlygate4sd3_1 hold569 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][9] ),
    .X(net1326));
 sg13g2_dlygate4sd3_1 hold570 (.A(_2537_),
    .X(net1327));
 sg13g2_dlygate4sd3_1 hold571 (.A(_0385_),
    .X(net1328));
 sg13g2_dlygate4sd3_1 hold572 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][4] ),
    .X(net1329));
 sg13g2_dlygate4sd3_1 hold573 (.A(_2833_),
    .X(net1330));
 sg13g2_dlygate4sd3_1 hold574 (.A(_0445_),
    .X(net1331));
 sg13g2_dlygate4sd3_1 hold575 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][6] ),
    .X(net1332));
 sg13g2_dlygate4sd3_1 hold576 (.A(_0153_),
    .X(net1333));
 sg13g2_dlygate4sd3_1 hold577 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][8] ),
    .X(net1334));
 sg13g2_dlygate4sd3_1 hold578 (.A(_2326_),
    .X(net1335));
 sg13g2_dlygate4sd3_1 hold579 (.A(_0346_),
    .X(net1336));
 sg13g2_dlygate4sd3_1 hold580 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][2] ),
    .X(net1337));
 sg13g2_dlygate4sd3_1 hold581 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][3] ),
    .X(net1338));
 sg13g2_dlygate4sd3_1 hold582 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][3] ),
    .X(net1339));
 sg13g2_dlygate4sd3_1 hold583 (.A(_0417_),
    .X(net1340));
 sg13g2_dlygate4sd3_1 hold584 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][11] ),
    .X(net1341));
 sg13g2_dlygate4sd3_1 hold585 (.A(_0222_),
    .X(net1342));
 sg13g2_dlygate4sd3_1 hold586 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[10] ),
    .X(net1343));
 sg13g2_dlygate4sd3_1 hold587 (.A(_2812_),
    .X(net1344));
 sg13g2_dlygate4sd3_1 hold588 (.A(_0438_),
    .X(net1345));
 sg13g2_dlygate4sd3_1 hold589 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][7] ),
    .X(net1346));
 sg13g2_dlygate4sd3_1 hold590 (.A(_2523_),
    .X(net1347));
 sg13g2_dlygate4sd3_1 hold591 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][4] ),
    .X(net1348));
 sg13g2_dlygate4sd3_1 hold592 (.A(_0380_),
    .X(net1349));
 sg13g2_dlygate4sd3_1 hold593 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][3] ),
    .X(net1350));
 sg13g2_dlygate4sd3_1 hold594 (.A(_1510_),
    .X(net1351));
 sg13g2_dlygate4sd3_1 hold595 (.A(_1511_),
    .X(net1352));
 sg13g2_dlygate4sd3_1 hold596 (.A(_0174_),
    .X(net1353));
 sg13g2_dlygate4sd3_1 hold597 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][6] ),
    .X(net1354));
 sg13g2_dlygate4sd3_1 hold598 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][2] ),
    .X(net1355));
 sg13g2_dlygate4sd3_1 hold599 (.A(_1127_),
    .X(net1356));
 sg13g2_dlygate4sd3_1 hold600 (.A(_0097_),
    .X(net1357));
 sg13g2_dlygate4sd3_1 hold601 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][4] ),
    .X(net1358));
 sg13g2_dlygate4sd3_1 hold602 (.A(_0331_),
    .X(net1359));
 sg13g2_dlygate4sd3_1 hold603 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][11] ),
    .X(net1360));
 sg13g2_dlygate4sd3_1 hold604 (.A(_1252_),
    .X(net1361));
 sg13g2_dlygate4sd3_1 hold605 (.A(_0119_),
    .X(net1362));
 sg13g2_dlygate4sd3_1 hold606 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][3] ),
    .X(net1363));
 sg13g2_dlygate4sd3_1 hold607 (.A(_1134_),
    .X(net1364));
 sg13g2_dlygate4sd3_1 hold608 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][1] ),
    .X(net1365));
 sg13g2_dlygate4sd3_1 hold609 (.A(_0199_),
    .X(net1366));
 sg13g2_dlygate4sd3_1 hold610 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[4][3] ),
    .X(net1367));
 sg13g2_dlygate4sd3_1 hold611 (.A(_0316_),
    .X(net1368));
 sg13g2_dlygate4sd3_1 hold612 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[2] ),
    .X(net1369));
 sg13g2_dlygate4sd3_1 hold613 (.A(_1362_),
    .X(net1370));
 sg13g2_dlygate4sd3_1 hold614 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][9] ),
    .X(net1371));
 sg13g2_dlygate4sd3_1 hold615 (.A(_2722_),
    .X(net1372));
 sg13g2_dlygate4sd3_1 hold616 (.A(_0424_),
    .X(net1373));
 sg13g2_dlygate4sd3_1 hold617 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][4] ),
    .X(net1374));
 sg13g2_dlygate4sd3_1 hold618 (.A(_1332_),
    .X(net1375));
 sg13g2_dlygate4sd3_1 hold619 (.A(_0137_),
    .X(net1376));
 sg13g2_dlygate4sd3_1 hold620 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[2] ),
    .X(net1377));
 sg13g2_dlygate4sd3_1 hold621 (.A(_0356_),
    .X(net1378));
 sg13g2_dlygate4sd3_1 hold622 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[4][2] ),
    .X(net1379));
 sg13g2_dlygate4sd3_1 hold623 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[5][4] ),
    .X(net1380));
 sg13g2_dlygate4sd3_1 hold624 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[3] ),
    .X(net1381));
 sg13g2_dlygate4sd3_1 hold625 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][2] ),
    .X(net1382));
 sg13g2_dlygate4sd3_1 hold626 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][3] ),
    .X(net1383));
 sg13g2_dlygate4sd3_1 hold627 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][3] ),
    .X(net1384));
 sg13g2_dlygate4sd3_1 hold628 (.A(_2290_),
    .X(net1385));
 sg13g2_dlygate4sd3_1 hold629 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][11] ),
    .X(net1386));
 sg13g2_dlygate4sd3_1 hold630 (.A(_0311_),
    .X(net1387));
 sg13g2_dlygate4sd3_1 hold631 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[3] ),
    .X(net1388));
 sg13g2_dlygate4sd3_1 hold632 (.A(_0320_),
    .X(net1389));
 sg13g2_dlygate4sd3_1 hold633 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][9] ),
    .X(net1390));
 sg13g2_dlygate4sd3_1 hold634 (.A(_0309_),
    .X(net1391));
 sg13g2_dlygate4sd3_1 hold635 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[1][9] ),
    .X(net1392));
 sg13g2_dlygate4sd3_1 hold636 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][2] ),
    .X(net1393));
 sg13g2_dlygate4sd3_1 hold637 (.A(_1897_),
    .X(net1394));
 sg13g2_dlygate4sd3_1 hold638 (.A(_0264_),
    .X(net1395));
 sg13g2_dlygate4sd3_1 hold639 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][5] ),
    .X(net1396));
 sg13g2_dlygate4sd3_1 hold640 (.A(_0241_),
    .X(net1397));
 sg13g2_dlygate4sd3_1 hold641 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][5] ),
    .X(net1398));
 sg13g2_dlygate4sd3_1 hold642 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][12] ),
    .X(net1399));
 sg13g2_dlygate4sd3_1 hold643 (.A(_0196_),
    .X(net1400));
 sg13g2_dlygate4sd3_1 hold644 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][7] ),
    .X(net1401));
 sg13g2_dlygate4sd3_1 hold645 (.A(_2317_),
    .X(net1402));
 sg13g2_dlygate4sd3_1 hold646 (.A(_0345_),
    .X(net1403));
 sg13g2_dlygate4sd3_1 hold647 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][5] ),
    .X(net1404));
 sg13g2_dlygate4sd3_1 hold648 (.A(_0113_),
    .X(net1405));
 sg13g2_dlygate4sd3_1 hold649 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[4] ),
    .X(net1406));
 sg13g2_dlygate4sd3_1 hold650 (.A(_0432_),
    .X(net1407));
 sg13g2_dlygate4sd3_1 hold651 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][12] ),
    .X(net1408));
 sg13g2_dlygate4sd3_1 hold652 (.A(_0274_),
    .X(net1409));
 sg13g2_dlygate4sd3_1 hold653 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][7] ),
    .X(net1410));
 sg13g2_dlygate4sd3_1 hold654 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][5] ),
    .X(net1411));
 sg13g2_dlygate4sd3_1 hold655 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][6] ),
    .X(net1412));
 sg13g2_dlygate4sd3_1 hold656 (.A(_2310_),
    .X(net1413));
 sg13g2_dlygate4sd3_1 hold657 (.A(_0344_),
    .X(net1414));
 sg13g2_dlygate4sd3_1 hold658 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][4] ),
    .X(net1415));
 sg13g2_dlygate4sd3_1 hold659 (.A(_0343_),
    .X(net1416));
 sg13g2_dlygate4sd3_1 hold660 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][5] ),
    .X(net1417));
 sg13g2_dlygate4sd3_1 hold661 (.A(_0305_),
    .X(net1418));
 sg13g2_dlygate4sd3_1 hold662 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[8][3] ),
    .X(net1419));
 sg13g2_dlygate4sd3_1 hold663 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[5] ),
    .X(net1420));
 sg13g2_dlygate4sd3_1 hold664 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][8] ),
    .X(net1421));
 sg13g2_dlygate4sd3_1 hold665 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][10] ),
    .X(net1422));
 sg13g2_dlygate4sd3_1 hold666 (.A(_2543_),
    .X(net1423));
 sg13g2_dlygate4sd3_1 hold667 (.A(_0386_),
    .X(net1424));
 sg13g2_dlygate4sd3_1 hold668 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[6] ),
    .X(net1425));
 sg13g2_dlygate4sd3_1 hold669 (.A(_2784_),
    .X(net1426));
 sg13g2_dlygate4sd3_1 hold670 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][1] ),
    .X(net1427));
 sg13g2_dlygate4sd3_1 hold671 (.A(_2477_),
    .X(net1428));
 sg13g2_dlygate4sd3_1 hold672 (.A(_0378_),
    .X(net1429));
 sg13g2_dlygate4sd3_1 hold673 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][7] ),
    .X(net1430));
 sg13g2_dlygate4sd3_1 hold674 (.A(_0243_),
    .X(net1431));
 sg13g2_dlygate4sd3_1 hold675 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][6] ),
    .X(net1432));
 sg13g2_dlygate4sd3_1 hold676 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][7] ),
    .X(net1433));
 sg13g2_dlygate4sd3_1 hold677 (.A(_1810_),
    .X(net1434));
 sg13g2_dlygate4sd3_1 hold678 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[6] ),
    .X(net1435));
 sg13g2_dlygate4sd3_1 hold679 (.A(_2606_),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold680 (.A(_0397_),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold681 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][2] ),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold682 (.A(_1574_),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold683 (.A(_0186_),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold684 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][4] ),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold685 (.A(_1406_),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold686 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[1] ),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold687 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][7] ),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold688 (.A(_0307_),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold689 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[3][2] ),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold690 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][3] ),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold691 (.A(_0214_),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold692 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[6] ),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold693 (.A(_2413_),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold694 (.A(_0360_),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold695 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][3] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold696 (.A(_0136_),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold697 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[4] ),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold698 (.A(_2593_),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold699 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[3] ),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold700 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[7] ),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold701 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][7] ),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold702 (.A(_1609_),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold703 (.A(_0192_),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold704 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][5] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold705 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][7] ),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold706 (.A(_1237_),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold707 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][2] ),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold708 (.A(_1786_),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold709 (.A(_0227_),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold710 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][10] ),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold711 (.A(_2339_),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold712 (.A(_0348_),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold713 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][2] ),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold714 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][6] ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold715 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[1] ),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold716 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[5][5] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold717 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][2] ),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold718 (.A(_2485_),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold719 (.A(_0379_),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold720 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][8] ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold721 (.A(_0155_),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold722 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][10] ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold723 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[7].y_shr[4] ),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold724 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][4] ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold725 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[3][9] ),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold726 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[6] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold727 (.A(_2220_),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold728 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][3] ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold729 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][11] ),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold730 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[3][8] ),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold731 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][2] ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold732 (.A(_1839_),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold733 (.A(_0238_),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold734 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[8] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold735 (.A(_0436_),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold736 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[9].y_shr[10] ),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold737 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][3] ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold738 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][6] ),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold739 (.A(_1599_),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold740 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][8] ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold741 (.A(_2716_),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold742 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[6][4] ),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold743 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][3] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold744 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][4] ),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold745 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[4] ),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold746 (.A(_0322_),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold747 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][9] ),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold748 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][4] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold749 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][6] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold750 (.A(_2256_),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold751 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[9] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold752 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[1] ),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold753 (.A(_2572_),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold754 (.A(_0392_),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold755 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][9] ),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold756 (.A(_0117_),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold757 (.A(\u_angle_cordic_12b_pmod.waveform_sel_reg[1] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold758 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][7] ),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold759 (.A(_1680_),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold760 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][2] ),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold761 (.A(_0302_),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold762 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[4] ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold763 (.A(_2406_),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold764 (.A(_0359_),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold765 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][6] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold766 (.A(_2694_),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold767 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][4] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold768 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[7][2] ),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold769 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[8][8] ),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold770 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][10] ),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold771 (.A(_1250_),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold772 (.A(_0118_),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold773 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[8] ),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold774 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[9] ),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold775 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][9] ),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold776 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][5] ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold777 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[8].y_shr[2] ),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold778 (.A(_1552_),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold779 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[7] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold780 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[7][7] ),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold781 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[1] ),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold782 (.A(_2012_),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold783 (.A(_0282_),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold784 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][6] ),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold785 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[0] ),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold786 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][4] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold787 (.A(_1799_),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold788 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[9][5] ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold789 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[3] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold790 (.A(_2761_),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold791 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][10] ),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold792 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[3].y_shr[7] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold793 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[8][5] ),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold794 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[5].y_shr[2] ),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold795 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[1].y_shr[1] ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold796 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][5] ),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold797 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[5] ),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold798 (.A(_0396_),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold799 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][2] ),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold800 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[1][10] ),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold801 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[5][8] ),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold802 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[3] ),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold803 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[10][6] ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold804 (.A(_0242_),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold805 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][8] ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold806 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.z[4][5] ),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold807 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][10] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold808 (.A(_1757_),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold809 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[4].y_shr[2] ),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold810 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][7] ),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold811 (.A(_1240_),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold812 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[9][12] ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold813 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[4][9] ),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold814 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[2].y_shr[7] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold815 (.A(_0383_),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold816 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.y[10][5] ),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold817 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[6][9] ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold818 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.x[2][8] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold819 (.A(\u_angle_cordic_12b_pmod.angle_cordic_12b.cordic.xyz[6].y_shr[3] ),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold820 (.A(\u_angle_cordic_12b_pmod.u_vga_top.v_cnt[0] ),
    .X(net1577));
 sg13g2_fill_1 FILLER_0_0 ();
 sg13g2_fill_2 FILLER_0_47 ();
 sg13g2_fill_2 FILLER_0_76 ();
 sg13g2_fill_1 FILLER_0_105 ();
 sg13g2_fill_2 FILLER_0_131 ();
 sg13g2_fill_1 FILLER_0_133 ();
 sg13g2_fill_2 FILLER_0_172 ();
 sg13g2_fill_1 FILLER_0_174 ();
 sg13g2_fill_2 FILLER_0_211 ();
 sg13g2_fill_1 FILLER_0_213 ();
 sg13g2_fill_2 FILLER_0_273 ();
 sg13g2_fill_1 FILLER_0_302 ();
 sg13g2_fill_2 FILLER_0_360 ();
 sg13g2_fill_2 FILLER_0_486 ();
 sg13g2_fill_1 FILLER_0_488 ();
 sg13g2_fill_2 FILLER_0_503 ();
 sg13g2_fill_2 FILLER_0_514 ();
 sg13g2_fill_2 FILLER_0_520 ();
 sg13g2_fill_1 FILLER_0_522 ();
 sg13g2_fill_1 FILLER_0_535 ();
 sg13g2_fill_2 FILLER_0_551 ();
 sg13g2_decap_8 FILLER_0_626 ();
 sg13g2_decap_8 FILLER_0_633 ();
 sg13g2_fill_2 FILLER_0_640 ();
 sg13g2_fill_1 FILLER_0_642 ();
 sg13g2_decap_8 FILLER_0_647 ();
 sg13g2_decap_8 FILLER_0_654 ();
 sg13g2_decap_8 FILLER_0_661 ();
 sg13g2_decap_8 FILLER_0_668 ();
 sg13g2_decap_8 FILLER_0_675 ();
 sg13g2_decap_8 FILLER_0_682 ();
 sg13g2_decap_8 FILLER_0_689 ();
 sg13g2_decap_8 FILLER_0_696 ();
 sg13g2_decap_8 FILLER_0_703 ();
 sg13g2_decap_8 FILLER_0_710 ();
 sg13g2_decap_8 FILLER_0_717 ();
 sg13g2_decap_8 FILLER_0_724 ();
 sg13g2_decap_8 FILLER_0_731 ();
 sg13g2_decap_8 FILLER_0_738 ();
 sg13g2_decap_8 FILLER_0_745 ();
 sg13g2_decap_8 FILLER_0_752 ();
 sg13g2_decap_8 FILLER_0_759 ();
 sg13g2_decap_8 FILLER_0_766 ();
 sg13g2_decap_8 FILLER_0_773 ();
 sg13g2_decap_8 FILLER_0_780 ();
 sg13g2_decap_8 FILLER_0_787 ();
 sg13g2_decap_8 FILLER_0_794 ();
 sg13g2_decap_8 FILLER_0_801 ();
 sg13g2_decap_8 FILLER_0_808 ();
 sg13g2_decap_8 FILLER_0_815 ();
 sg13g2_decap_8 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_0_829 ();
 sg13g2_decap_8 FILLER_0_836 ();
 sg13g2_decap_8 FILLER_0_843 ();
 sg13g2_decap_8 FILLER_0_850 ();
 sg13g2_decap_8 FILLER_0_857 ();
 sg13g2_decap_8 FILLER_0_864 ();
 sg13g2_decap_8 FILLER_0_871 ();
 sg13g2_decap_8 FILLER_0_878 ();
 sg13g2_decap_8 FILLER_0_885 ();
 sg13g2_decap_8 FILLER_0_892 ();
 sg13g2_decap_8 FILLER_0_899 ();
 sg13g2_decap_8 FILLER_0_906 ();
 sg13g2_decap_8 FILLER_0_913 ();
 sg13g2_decap_8 FILLER_0_920 ();
 sg13g2_decap_8 FILLER_0_927 ();
 sg13g2_decap_8 FILLER_0_934 ();
 sg13g2_decap_8 FILLER_0_941 ();
 sg13g2_decap_8 FILLER_0_948 ();
 sg13g2_decap_8 FILLER_0_955 ();
 sg13g2_decap_8 FILLER_0_962 ();
 sg13g2_decap_8 FILLER_0_969 ();
 sg13g2_decap_8 FILLER_0_976 ();
 sg13g2_decap_8 FILLER_0_983 ();
 sg13g2_decap_8 FILLER_0_990 ();
 sg13g2_decap_8 FILLER_0_997 ();
 sg13g2_decap_8 FILLER_0_1004 ();
 sg13g2_decap_8 FILLER_0_1011 ();
 sg13g2_decap_8 FILLER_0_1018 ();
 sg13g2_decap_4 FILLER_0_1025 ();
 sg13g2_fill_2 FILLER_1_0 ();
 sg13g2_fill_1 FILLER_1_183 ();
 sg13g2_fill_2 FILLER_1_220 ();
 sg13g2_fill_1 FILLER_1_222 ();
 sg13g2_fill_2 FILLER_1_260 ();
 sg13g2_fill_2 FILLER_1_279 ();
 sg13g2_fill_1 FILLER_1_281 ();
 sg13g2_fill_2 FILLER_1_295 ();
 sg13g2_fill_2 FILLER_1_318 ();
 sg13g2_fill_1 FILLER_1_329 ();
 sg13g2_fill_1 FILLER_1_358 ();
 sg13g2_fill_1 FILLER_1_372 ();
 sg13g2_fill_2 FILLER_1_541 ();
 sg13g2_fill_1 FILLER_1_561 ();
 sg13g2_fill_1 FILLER_1_626 ();
 sg13g2_fill_1 FILLER_1_636 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_decap_8 FILLER_1_875 ();
 sg13g2_decap_8 FILLER_1_882 ();
 sg13g2_decap_8 FILLER_1_889 ();
 sg13g2_decap_8 FILLER_1_896 ();
 sg13g2_decap_8 FILLER_1_903 ();
 sg13g2_decap_8 FILLER_1_910 ();
 sg13g2_decap_8 FILLER_1_917 ();
 sg13g2_decap_8 FILLER_1_924 ();
 sg13g2_decap_8 FILLER_1_931 ();
 sg13g2_decap_8 FILLER_1_938 ();
 sg13g2_decap_8 FILLER_1_945 ();
 sg13g2_decap_8 FILLER_1_952 ();
 sg13g2_decap_8 FILLER_1_959 ();
 sg13g2_decap_8 FILLER_1_966 ();
 sg13g2_decap_8 FILLER_1_973 ();
 sg13g2_decap_8 FILLER_1_980 ();
 sg13g2_decap_8 FILLER_1_987 ();
 sg13g2_decap_8 FILLER_1_994 ();
 sg13g2_decap_8 FILLER_1_1001 ();
 sg13g2_decap_8 FILLER_1_1008 ();
 sg13g2_decap_8 FILLER_1_1015 ();
 sg13g2_decap_8 FILLER_1_1022 ();
 sg13g2_fill_2 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_102 ();
 sg13g2_fill_2 FILLER_2_144 ();
 sg13g2_fill_2 FILLER_2_192 ();
 sg13g2_fill_2 FILLER_2_291 ();
 sg13g2_fill_2 FILLER_2_376 ();
 sg13g2_fill_1 FILLER_2_387 ();
 sg13g2_fill_1 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_421 ();
 sg13g2_fill_2 FILLER_2_464 ();
 sg13g2_fill_1 FILLER_2_466 ();
 sg13g2_fill_1 FILLER_2_514 ();
 sg13g2_fill_1 FILLER_2_525 ();
 sg13g2_fill_2 FILLER_2_545 ();
 sg13g2_fill_1 FILLER_2_578 ();
 sg13g2_fill_1 FILLER_2_610 ();
 sg13g2_decap_8 FILLER_2_669 ();
 sg13g2_decap_8 FILLER_2_676 ();
 sg13g2_decap_8 FILLER_2_683 ();
 sg13g2_decap_8 FILLER_2_690 ();
 sg13g2_decap_8 FILLER_2_697 ();
 sg13g2_decap_8 FILLER_2_704 ();
 sg13g2_decap_8 FILLER_2_711 ();
 sg13g2_decap_8 FILLER_2_718 ();
 sg13g2_decap_8 FILLER_2_725 ();
 sg13g2_decap_8 FILLER_2_732 ();
 sg13g2_decap_8 FILLER_2_739 ();
 sg13g2_decap_8 FILLER_2_746 ();
 sg13g2_decap_8 FILLER_2_753 ();
 sg13g2_decap_8 FILLER_2_760 ();
 sg13g2_decap_8 FILLER_2_767 ();
 sg13g2_decap_8 FILLER_2_774 ();
 sg13g2_decap_8 FILLER_2_781 ();
 sg13g2_decap_8 FILLER_2_788 ();
 sg13g2_decap_8 FILLER_2_795 ();
 sg13g2_decap_8 FILLER_2_802 ();
 sg13g2_decap_8 FILLER_2_809 ();
 sg13g2_decap_8 FILLER_2_816 ();
 sg13g2_decap_8 FILLER_2_823 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_844 ();
 sg13g2_decap_8 FILLER_2_851 ();
 sg13g2_decap_8 FILLER_2_858 ();
 sg13g2_decap_8 FILLER_2_865 ();
 sg13g2_decap_8 FILLER_2_872 ();
 sg13g2_decap_8 FILLER_2_879 ();
 sg13g2_decap_8 FILLER_2_886 ();
 sg13g2_decap_8 FILLER_2_893 ();
 sg13g2_decap_8 FILLER_2_900 ();
 sg13g2_decap_8 FILLER_2_907 ();
 sg13g2_decap_8 FILLER_2_914 ();
 sg13g2_decap_8 FILLER_2_921 ();
 sg13g2_decap_8 FILLER_2_928 ();
 sg13g2_decap_8 FILLER_2_935 ();
 sg13g2_decap_8 FILLER_2_942 ();
 sg13g2_decap_8 FILLER_2_949 ();
 sg13g2_decap_8 FILLER_2_956 ();
 sg13g2_decap_8 FILLER_2_963 ();
 sg13g2_decap_8 FILLER_2_970 ();
 sg13g2_decap_8 FILLER_2_977 ();
 sg13g2_decap_8 FILLER_2_984 ();
 sg13g2_decap_8 FILLER_2_991 ();
 sg13g2_decap_8 FILLER_2_998 ();
 sg13g2_decap_8 FILLER_2_1005 ();
 sg13g2_decap_8 FILLER_2_1012 ();
 sg13g2_decap_8 FILLER_2_1019 ();
 sg13g2_fill_2 FILLER_2_1026 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_fill_2 FILLER_3_83 ();
 sg13g2_fill_1 FILLER_3_112 ();
 sg13g2_fill_2 FILLER_3_256 ();
 sg13g2_fill_1 FILLER_3_258 ();
 sg13g2_fill_1 FILLER_3_336 ();
 sg13g2_fill_1 FILLER_3_391 ();
 sg13g2_fill_1 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_451 ();
 sg13g2_fill_2 FILLER_3_508 ();
 sg13g2_fill_1 FILLER_3_515 ();
 sg13g2_fill_2 FILLER_3_543 ();
 sg13g2_fill_2 FILLER_3_558 ();
 sg13g2_fill_1 FILLER_3_591 ();
 sg13g2_fill_1 FILLER_3_601 ();
 sg13g2_fill_1 FILLER_3_611 ();
 sg13g2_fill_2 FILLER_3_640 ();
 sg13g2_decap_8 FILLER_3_682 ();
 sg13g2_decap_8 FILLER_3_689 ();
 sg13g2_decap_8 FILLER_3_696 ();
 sg13g2_decap_8 FILLER_3_703 ();
 sg13g2_decap_8 FILLER_3_710 ();
 sg13g2_decap_8 FILLER_3_717 ();
 sg13g2_decap_8 FILLER_3_724 ();
 sg13g2_decap_8 FILLER_3_731 ();
 sg13g2_decap_8 FILLER_3_738 ();
 sg13g2_decap_8 FILLER_3_745 ();
 sg13g2_decap_8 FILLER_3_752 ();
 sg13g2_decap_8 FILLER_3_759 ();
 sg13g2_decap_8 FILLER_3_766 ();
 sg13g2_decap_8 FILLER_3_773 ();
 sg13g2_decap_8 FILLER_3_780 ();
 sg13g2_decap_8 FILLER_3_787 ();
 sg13g2_decap_8 FILLER_3_794 ();
 sg13g2_decap_8 FILLER_3_801 ();
 sg13g2_decap_8 FILLER_3_808 ();
 sg13g2_decap_8 FILLER_3_815 ();
 sg13g2_decap_8 FILLER_3_822 ();
 sg13g2_decap_8 FILLER_3_829 ();
 sg13g2_decap_8 FILLER_3_836 ();
 sg13g2_decap_8 FILLER_3_843 ();
 sg13g2_decap_8 FILLER_3_850 ();
 sg13g2_decap_8 FILLER_3_857 ();
 sg13g2_decap_8 FILLER_3_864 ();
 sg13g2_decap_8 FILLER_3_871 ();
 sg13g2_decap_8 FILLER_3_878 ();
 sg13g2_decap_8 FILLER_3_885 ();
 sg13g2_decap_8 FILLER_3_892 ();
 sg13g2_decap_8 FILLER_3_899 ();
 sg13g2_decap_8 FILLER_3_906 ();
 sg13g2_decap_8 FILLER_3_913 ();
 sg13g2_decap_8 FILLER_3_920 ();
 sg13g2_decap_8 FILLER_3_927 ();
 sg13g2_decap_8 FILLER_3_934 ();
 sg13g2_decap_8 FILLER_3_941 ();
 sg13g2_decap_8 FILLER_3_948 ();
 sg13g2_decap_8 FILLER_3_955 ();
 sg13g2_decap_8 FILLER_3_962 ();
 sg13g2_decap_8 FILLER_3_969 ();
 sg13g2_decap_8 FILLER_3_976 ();
 sg13g2_decap_8 FILLER_3_983 ();
 sg13g2_decap_8 FILLER_3_990 ();
 sg13g2_decap_8 FILLER_3_997 ();
 sg13g2_decap_8 FILLER_3_1004 ();
 sg13g2_decap_8 FILLER_3_1011 ();
 sg13g2_decap_8 FILLER_3_1018 ();
 sg13g2_decap_4 FILLER_3_1025 ();
 sg13g2_fill_2 FILLER_4_32 ();
 sg13g2_fill_2 FILLER_4_153 ();
 sg13g2_fill_1 FILLER_4_155 ();
 sg13g2_fill_1 FILLER_4_184 ();
 sg13g2_fill_2 FILLER_4_213 ();
 sg13g2_fill_1 FILLER_4_215 ();
 sg13g2_fill_2 FILLER_4_265 ();
 sg13g2_fill_2 FILLER_4_282 ();
 sg13g2_fill_1 FILLER_4_284 ();
 sg13g2_fill_2 FILLER_4_382 ();
 sg13g2_fill_2 FILLER_4_397 ();
 sg13g2_fill_2 FILLER_4_528 ();
 sg13g2_fill_2 FILLER_4_545 ();
 sg13g2_fill_1 FILLER_4_547 ();
 sg13g2_fill_1 FILLER_4_645 ();
 sg13g2_decap_8 FILLER_4_685 ();
 sg13g2_decap_8 FILLER_4_692 ();
 sg13g2_decap_8 FILLER_4_699 ();
 sg13g2_decap_8 FILLER_4_706 ();
 sg13g2_decap_8 FILLER_4_713 ();
 sg13g2_decap_8 FILLER_4_720 ();
 sg13g2_decap_8 FILLER_4_727 ();
 sg13g2_decap_8 FILLER_4_734 ();
 sg13g2_decap_8 FILLER_4_741 ();
 sg13g2_decap_8 FILLER_4_748 ();
 sg13g2_decap_8 FILLER_4_755 ();
 sg13g2_decap_8 FILLER_4_762 ();
 sg13g2_decap_8 FILLER_4_769 ();
 sg13g2_decap_8 FILLER_4_776 ();
 sg13g2_decap_8 FILLER_4_783 ();
 sg13g2_decap_8 FILLER_4_790 ();
 sg13g2_decap_8 FILLER_4_797 ();
 sg13g2_decap_8 FILLER_4_804 ();
 sg13g2_decap_8 FILLER_4_811 ();
 sg13g2_decap_8 FILLER_4_818 ();
 sg13g2_decap_8 FILLER_4_825 ();
 sg13g2_decap_8 FILLER_4_832 ();
 sg13g2_decap_8 FILLER_4_839 ();
 sg13g2_decap_8 FILLER_4_846 ();
 sg13g2_decap_8 FILLER_4_853 ();
 sg13g2_decap_8 FILLER_4_860 ();
 sg13g2_decap_8 FILLER_4_867 ();
 sg13g2_decap_8 FILLER_4_874 ();
 sg13g2_decap_8 FILLER_4_881 ();
 sg13g2_decap_8 FILLER_4_888 ();
 sg13g2_decap_8 FILLER_4_895 ();
 sg13g2_decap_8 FILLER_4_902 ();
 sg13g2_decap_8 FILLER_4_909 ();
 sg13g2_decap_8 FILLER_4_916 ();
 sg13g2_decap_8 FILLER_4_923 ();
 sg13g2_decap_8 FILLER_4_930 ();
 sg13g2_decap_8 FILLER_4_937 ();
 sg13g2_decap_8 FILLER_4_944 ();
 sg13g2_decap_8 FILLER_4_951 ();
 sg13g2_decap_8 FILLER_4_958 ();
 sg13g2_decap_8 FILLER_4_965 ();
 sg13g2_decap_8 FILLER_4_972 ();
 sg13g2_decap_8 FILLER_4_979 ();
 sg13g2_decap_8 FILLER_4_986 ();
 sg13g2_decap_8 FILLER_4_993 ();
 sg13g2_decap_8 FILLER_4_1000 ();
 sg13g2_decap_8 FILLER_4_1007 ();
 sg13g2_decap_8 FILLER_4_1014 ();
 sg13g2_decap_8 FILLER_4_1021 ();
 sg13g2_fill_1 FILLER_4_1028 ();
 sg13g2_fill_1 FILLER_5_57 ();
 sg13g2_fill_2 FILLER_5_63 ();
 sg13g2_fill_2 FILLER_5_100 ();
 sg13g2_fill_2 FILLER_5_134 ();
 sg13g2_fill_2 FILLER_5_164 ();
 sg13g2_fill_2 FILLER_5_190 ();
 sg13g2_fill_2 FILLER_5_201 ();
 sg13g2_fill_1 FILLER_5_250 ();
 sg13g2_fill_1 FILLER_5_265 ();
 sg13g2_fill_1 FILLER_5_271 ();
 sg13g2_fill_1 FILLER_5_323 ();
 sg13g2_fill_2 FILLER_5_377 ();
 sg13g2_fill_1 FILLER_5_435 ();
 sg13g2_fill_2 FILLER_5_469 ();
 sg13g2_fill_1 FILLER_5_502 ();
 sg13g2_fill_2 FILLER_5_566 ();
 sg13g2_fill_1 FILLER_5_568 ();
 sg13g2_fill_1 FILLER_5_623 ();
 sg13g2_fill_2 FILLER_5_666 ();
 sg13g2_fill_1 FILLER_5_668 ();
 sg13g2_decap_8 FILLER_5_709 ();
 sg13g2_decap_8 FILLER_5_716 ();
 sg13g2_decap_8 FILLER_5_723 ();
 sg13g2_decap_8 FILLER_5_730 ();
 sg13g2_decap_8 FILLER_5_737 ();
 sg13g2_decap_8 FILLER_5_744 ();
 sg13g2_decap_8 FILLER_5_751 ();
 sg13g2_decap_8 FILLER_5_758 ();
 sg13g2_decap_8 FILLER_5_765 ();
 sg13g2_decap_8 FILLER_5_772 ();
 sg13g2_decap_8 FILLER_5_779 ();
 sg13g2_decap_8 FILLER_5_786 ();
 sg13g2_decap_8 FILLER_5_793 ();
 sg13g2_decap_8 FILLER_5_800 ();
 sg13g2_decap_8 FILLER_5_807 ();
 sg13g2_decap_8 FILLER_5_814 ();
 sg13g2_decap_8 FILLER_5_821 ();
 sg13g2_decap_8 FILLER_5_828 ();
 sg13g2_decap_8 FILLER_5_835 ();
 sg13g2_decap_8 FILLER_5_842 ();
 sg13g2_decap_8 FILLER_5_849 ();
 sg13g2_decap_8 FILLER_5_856 ();
 sg13g2_decap_8 FILLER_5_863 ();
 sg13g2_decap_8 FILLER_5_870 ();
 sg13g2_decap_8 FILLER_5_877 ();
 sg13g2_decap_8 FILLER_5_884 ();
 sg13g2_decap_8 FILLER_5_891 ();
 sg13g2_decap_8 FILLER_5_898 ();
 sg13g2_decap_8 FILLER_5_905 ();
 sg13g2_decap_8 FILLER_5_912 ();
 sg13g2_decap_8 FILLER_5_919 ();
 sg13g2_decap_8 FILLER_5_926 ();
 sg13g2_decap_8 FILLER_5_933 ();
 sg13g2_decap_8 FILLER_5_940 ();
 sg13g2_decap_8 FILLER_5_947 ();
 sg13g2_decap_8 FILLER_5_954 ();
 sg13g2_decap_8 FILLER_5_961 ();
 sg13g2_decap_8 FILLER_5_968 ();
 sg13g2_decap_8 FILLER_5_975 ();
 sg13g2_decap_8 FILLER_5_982 ();
 sg13g2_decap_8 FILLER_5_989 ();
 sg13g2_decap_8 FILLER_5_996 ();
 sg13g2_decap_8 FILLER_5_1003 ();
 sg13g2_decap_8 FILLER_5_1010 ();
 sg13g2_decap_8 FILLER_5_1017 ();
 sg13g2_decap_4 FILLER_5_1024 ();
 sg13g2_fill_1 FILLER_5_1028 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_38 ();
 sg13g2_fill_1 FILLER_6_123 ();
 sg13g2_fill_1 FILLER_6_211 ();
 sg13g2_fill_1 FILLER_6_247 ();
 sg13g2_fill_1 FILLER_6_377 ();
 sg13g2_fill_1 FILLER_6_397 ();
 sg13g2_fill_1 FILLER_6_413 ();
 sg13g2_fill_2 FILLER_6_453 ();
 sg13g2_fill_2 FILLER_6_500 ();
 sg13g2_fill_1 FILLER_6_540 ();
 sg13g2_fill_2 FILLER_6_621 ();
 sg13g2_fill_2 FILLER_6_632 ();
 sg13g2_fill_1 FILLER_6_634 ();
 sg13g2_decap_4 FILLER_6_701 ();
 sg13g2_decap_8 FILLER_6_709 ();
 sg13g2_decap_8 FILLER_6_720 ();
 sg13g2_decap_8 FILLER_6_727 ();
 sg13g2_decap_8 FILLER_6_734 ();
 sg13g2_decap_8 FILLER_6_741 ();
 sg13g2_decap_8 FILLER_6_748 ();
 sg13g2_decap_8 FILLER_6_755 ();
 sg13g2_decap_8 FILLER_6_762 ();
 sg13g2_decap_8 FILLER_6_769 ();
 sg13g2_decap_8 FILLER_6_776 ();
 sg13g2_decap_8 FILLER_6_783 ();
 sg13g2_decap_8 FILLER_6_790 ();
 sg13g2_decap_8 FILLER_6_797 ();
 sg13g2_decap_8 FILLER_6_804 ();
 sg13g2_decap_8 FILLER_6_811 ();
 sg13g2_decap_8 FILLER_6_818 ();
 sg13g2_decap_8 FILLER_6_825 ();
 sg13g2_decap_8 FILLER_6_832 ();
 sg13g2_decap_8 FILLER_6_839 ();
 sg13g2_decap_8 FILLER_6_846 ();
 sg13g2_decap_8 FILLER_6_853 ();
 sg13g2_decap_8 FILLER_6_860 ();
 sg13g2_decap_8 FILLER_6_867 ();
 sg13g2_decap_8 FILLER_6_874 ();
 sg13g2_decap_8 FILLER_6_881 ();
 sg13g2_decap_8 FILLER_6_888 ();
 sg13g2_decap_8 FILLER_6_895 ();
 sg13g2_decap_8 FILLER_6_902 ();
 sg13g2_decap_8 FILLER_6_909 ();
 sg13g2_decap_8 FILLER_6_916 ();
 sg13g2_decap_8 FILLER_6_923 ();
 sg13g2_decap_8 FILLER_6_930 ();
 sg13g2_decap_8 FILLER_6_937 ();
 sg13g2_decap_8 FILLER_6_944 ();
 sg13g2_decap_8 FILLER_6_951 ();
 sg13g2_decap_8 FILLER_6_958 ();
 sg13g2_decap_8 FILLER_6_965 ();
 sg13g2_decap_8 FILLER_6_972 ();
 sg13g2_decap_8 FILLER_6_979 ();
 sg13g2_decap_8 FILLER_6_986 ();
 sg13g2_decap_8 FILLER_6_993 ();
 sg13g2_decap_8 FILLER_6_1000 ();
 sg13g2_decap_8 FILLER_6_1007 ();
 sg13g2_decap_8 FILLER_6_1014 ();
 sg13g2_decap_8 FILLER_6_1021 ();
 sg13g2_fill_1 FILLER_6_1028 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_51 ();
 sg13g2_fill_1 FILLER_7_108 ();
 sg13g2_fill_1 FILLER_7_205 ();
 sg13g2_fill_1 FILLER_7_282 ();
 sg13g2_fill_1 FILLER_7_293 ();
 sg13g2_fill_2 FILLER_7_321 ();
 sg13g2_fill_1 FILLER_7_323 ();
 sg13g2_fill_1 FILLER_7_351 ();
 sg13g2_fill_1 FILLER_7_371 ();
 sg13g2_fill_1 FILLER_7_405 ();
 sg13g2_fill_1 FILLER_7_415 ();
 sg13g2_fill_1 FILLER_7_434 ();
 sg13g2_fill_1 FILLER_7_462 ();
 sg13g2_fill_1 FILLER_7_467 ();
 sg13g2_fill_2 FILLER_7_495 ();
 sg13g2_fill_1 FILLER_7_527 ();
 sg13g2_fill_1 FILLER_7_563 ();
 sg13g2_fill_2 FILLER_7_611 ();
 sg13g2_fill_2 FILLER_7_621 ();
 sg13g2_fill_1 FILLER_7_623 ();
 sg13g2_fill_1 FILLER_7_647 ();
 sg13g2_fill_2 FILLER_7_706 ();
 sg13g2_fill_2 FILLER_7_725 ();
 sg13g2_fill_2 FILLER_7_735 ();
 sg13g2_fill_1 FILLER_7_737 ();
 sg13g2_decap_8 FILLER_7_746 ();
 sg13g2_decap_8 FILLER_7_753 ();
 sg13g2_decap_8 FILLER_7_760 ();
 sg13g2_decap_4 FILLER_7_767 ();
 sg13g2_fill_2 FILLER_7_775 ();
 sg13g2_decap_4 FILLER_7_781 ();
 sg13g2_fill_2 FILLER_7_785 ();
 sg13g2_decap_8 FILLER_7_799 ();
 sg13g2_decap_8 FILLER_7_806 ();
 sg13g2_decap_8 FILLER_7_813 ();
 sg13g2_decap_8 FILLER_7_820 ();
 sg13g2_decap_8 FILLER_7_827 ();
 sg13g2_decap_8 FILLER_7_834 ();
 sg13g2_decap_8 FILLER_7_841 ();
 sg13g2_decap_8 FILLER_7_848 ();
 sg13g2_decap_8 FILLER_7_855 ();
 sg13g2_decap_8 FILLER_7_862 ();
 sg13g2_decap_8 FILLER_7_869 ();
 sg13g2_decap_8 FILLER_7_876 ();
 sg13g2_decap_8 FILLER_7_883 ();
 sg13g2_decap_8 FILLER_7_890 ();
 sg13g2_decap_8 FILLER_7_897 ();
 sg13g2_decap_8 FILLER_7_904 ();
 sg13g2_decap_8 FILLER_7_911 ();
 sg13g2_decap_8 FILLER_7_918 ();
 sg13g2_decap_8 FILLER_7_925 ();
 sg13g2_decap_8 FILLER_7_932 ();
 sg13g2_decap_8 FILLER_7_939 ();
 sg13g2_decap_8 FILLER_7_946 ();
 sg13g2_decap_8 FILLER_7_953 ();
 sg13g2_decap_8 FILLER_7_960 ();
 sg13g2_decap_8 FILLER_7_967 ();
 sg13g2_decap_8 FILLER_7_974 ();
 sg13g2_decap_8 FILLER_7_981 ();
 sg13g2_decap_8 FILLER_7_988 ();
 sg13g2_decap_8 FILLER_7_995 ();
 sg13g2_decap_8 FILLER_7_1002 ();
 sg13g2_decap_8 FILLER_7_1009 ();
 sg13g2_decap_8 FILLER_7_1016 ();
 sg13g2_decap_4 FILLER_7_1023 ();
 sg13g2_fill_2 FILLER_7_1027 ();
 sg13g2_fill_2 FILLER_8_47 ();
 sg13g2_fill_1 FILLER_8_54 ();
 sg13g2_fill_1 FILLER_8_165 ();
 sg13g2_fill_2 FILLER_8_203 ();
 sg13g2_fill_1 FILLER_8_205 ();
 sg13g2_fill_2 FILLER_8_219 ();
 sg13g2_fill_1 FILLER_8_221 ();
 sg13g2_fill_1 FILLER_8_287 ();
 sg13g2_fill_1 FILLER_8_328 ();
 sg13g2_fill_2 FILLER_8_373 ();
 sg13g2_fill_1 FILLER_8_449 ();
 sg13g2_fill_1 FILLER_8_481 ();
 sg13g2_fill_1 FILLER_8_502 ();
 sg13g2_fill_1 FILLER_8_508 ();
 sg13g2_fill_2 FILLER_8_589 ();
 sg13g2_fill_2 FILLER_8_613 ();
 sg13g2_fill_1 FILLER_8_671 ();
 sg13g2_fill_2 FILLER_8_681 ();
 sg13g2_fill_2 FILLER_8_697 ();
 sg13g2_fill_1 FILLER_8_699 ();
 sg13g2_fill_1 FILLER_8_758 ();
 sg13g2_fill_2 FILLER_8_793 ();
 sg13g2_fill_1 FILLER_8_795 ();
 sg13g2_fill_1 FILLER_8_805 ();
 sg13g2_decap_4 FILLER_8_811 ();
 sg13g2_fill_1 FILLER_8_815 ();
 sg13g2_decap_8 FILLER_8_825 ();
 sg13g2_decap_8 FILLER_8_832 ();
 sg13g2_decap_8 FILLER_8_839 ();
 sg13g2_decap_8 FILLER_8_846 ();
 sg13g2_decap_8 FILLER_8_853 ();
 sg13g2_decap_8 FILLER_8_860 ();
 sg13g2_decap_8 FILLER_8_867 ();
 sg13g2_decap_8 FILLER_8_874 ();
 sg13g2_decap_8 FILLER_8_881 ();
 sg13g2_decap_8 FILLER_8_888 ();
 sg13g2_decap_8 FILLER_8_895 ();
 sg13g2_decap_8 FILLER_8_902 ();
 sg13g2_decap_8 FILLER_8_909 ();
 sg13g2_decap_8 FILLER_8_916 ();
 sg13g2_decap_8 FILLER_8_923 ();
 sg13g2_decap_8 FILLER_8_930 ();
 sg13g2_decap_8 FILLER_8_937 ();
 sg13g2_decap_8 FILLER_8_944 ();
 sg13g2_decap_8 FILLER_8_951 ();
 sg13g2_decap_8 FILLER_8_958 ();
 sg13g2_decap_8 FILLER_8_965 ();
 sg13g2_decap_8 FILLER_8_972 ();
 sg13g2_decap_8 FILLER_8_979 ();
 sg13g2_decap_8 FILLER_8_986 ();
 sg13g2_decap_8 FILLER_8_993 ();
 sg13g2_decap_8 FILLER_8_1000 ();
 sg13g2_decap_8 FILLER_8_1007 ();
 sg13g2_decap_8 FILLER_8_1014 ();
 sg13g2_decap_8 FILLER_8_1021 ();
 sg13g2_fill_1 FILLER_8_1028 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_90 ();
 sg13g2_fill_2 FILLER_9_140 ();
 sg13g2_fill_1 FILLER_9_142 ();
 sg13g2_fill_1 FILLER_9_179 ();
 sg13g2_fill_2 FILLER_9_349 ();
 sg13g2_fill_2 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_421 ();
 sg13g2_fill_1 FILLER_9_423 ();
 sg13g2_fill_2 FILLER_9_470 ();
 sg13g2_fill_1 FILLER_9_472 ();
 sg13g2_fill_1 FILLER_9_511 ();
 sg13g2_fill_2 FILLER_9_520 ();
 sg13g2_fill_2 FILLER_9_535 ();
 sg13g2_fill_1 FILLER_9_556 ();
 sg13g2_fill_2 FILLER_9_566 ();
 sg13g2_fill_2 FILLER_9_659 ();
 sg13g2_fill_2 FILLER_9_743 ();
 sg13g2_fill_1 FILLER_9_745 ();
 sg13g2_fill_2 FILLER_9_786 ();
 sg13g2_fill_1 FILLER_9_788 ();
 sg13g2_decap_8 FILLER_9_841 ();
 sg13g2_decap_8 FILLER_9_848 ();
 sg13g2_decap_8 FILLER_9_855 ();
 sg13g2_decap_8 FILLER_9_862 ();
 sg13g2_decap_8 FILLER_9_869 ();
 sg13g2_decap_8 FILLER_9_876 ();
 sg13g2_decap_8 FILLER_9_883 ();
 sg13g2_decap_8 FILLER_9_890 ();
 sg13g2_decap_8 FILLER_9_897 ();
 sg13g2_decap_8 FILLER_9_904 ();
 sg13g2_decap_8 FILLER_9_911 ();
 sg13g2_decap_8 FILLER_9_918 ();
 sg13g2_decap_8 FILLER_9_925 ();
 sg13g2_decap_8 FILLER_9_932 ();
 sg13g2_decap_8 FILLER_9_939 ();
 sg13g2_decap_8 FILLER_9_946 ();
 sg13g2_decap_8 FILLER_9_953 ();
 sg13g2_decap_8 FILLER_9_960 ();
 sg13g2_decap_8 FILLER_9_967 ();
 sg13g2_decap_8 FILLER_9_974 ();
 sg13g2_decap_8 FILLER_9_981 ();
 sg13g2_decap_8 FILLER_9_988 ();
 sg13g2_decap_8 FILLER_9_995 ();
 sg13g2_decap_8 FILLER_9_1002 ();
 sg13g2_decap_8 FILLER_9_1009 ();
 sg13g2_decap_8 FILLER_9_1016 ();
 sg13g2_decap_4 FILLER_9_1023 ();
 sg13g2_fill_2 FILLER_9_1027 ();
 sg13g2_fill_2 FILLER_10_36 ();
 sg13g2_fill_1 FILLER_10_116 ();
 sg13g2_fill_2 FILLER_10_130 ();
 sg13g2_fill_2 FILLER_10_202 ();
 sg13g2_fill_1 FILLER_10_204 ();
 sg13g2_fill_2 FILLER_10_297 ();
 sg13g2_fill_1 FILLER_10_436 ();
 sg13g2_fill_2 FILLER_10_485 ();
 sg13g2_fill_1 FILLER_10_519 ();
 sg13g2_fill_1 FILLER_10_602 ();
 sg13g2_fill_1 FILLER_10_653 ();
 sg13g2_fill_1 FILLER_10_667 ();
 sg13g2_fill_2 FILLER_10_692 ();
 sg13g2_fill_2 FILLER_10_720 ();
 sg13g2_fill_2 FILLER_10_794 ();
 sg13g2_fill_1 FILLER_10_796 ();
 sg13g2_decap_8 FILLER_10_852 ();
 sg13g2_decap_8 FILLER_10_859 ();
 sg13g2_decap_8 FILLER_10_866 ();
 sg13g2_decap_8 FILLER_10_873 ();
 sg13g2_decap_8 FILLER_10_880 ();
 sg13g2_decap_8 FILLER_10_887 ();
 sg13g2_decap_8 FILLER_10_894 ();
 sg13g2_decap_8 FILLER_10_901 ();
 sg13g2_decap_8 FILLER_10_908 ();
 sg13g2_decap_8 FILLER_10_915 ();
 sg13g2_decap_8 FILLER_10_922 ();
 sg13g2_decap_8 FILLER_10_929 ();
 sg13g2_decap_8 FILLER_10_936 ();
 sg13g2_decap_8 FILLER_10_943 ();
 sg13g2_decap_8 FILLER_10_950 ();
 sg13g2_decap_8 FILLER_10_957 ();
 sg13g2_decap_8 FILLER_10_964 ();
 sg13g2_decap_8 FILLER_10_971 ();
 sg13g2_decap_8 FILLER_10_978 ();
 sg13g2_decap_8 FILLER_10_985 ();
 sg13g2_decap_8 FILLER_10_992 ();
 sg13g2_decap_8 FILLER_10_999 ();
 sg13g2_decap_8 FILLER_10_1006 ();
 sg13g2_decap_8 FILLER_10_1013 ();
 sg13g2_decap_8 FILLER_10_1020 ();
 sg13g2_fill_2 FILLER_10_1027 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_2 ();
 sg13g2_fill_2 FILLER_11_62 ();
 sg13g2_fill_1 FILLER_11_64 ();
 sg13g2_fill_1 FILLER_11_84 ();
 sg13g2_fill_2 FILLER_11_113 ();
 sg13g2_fill_1 FILLER_11_143 ();
 sg13g2_fill_1 FILLER_11_153 ();
 sg13g2_fill_1 FILLER_11_217 ();
 sg13g2_fill_1 FILLER_11_280 ();
 sg13g2_fill_1 FILLER_11_338 ();
 sg13g2_fill_1 FILLER_11_413 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_fill_2 FILLER_11_519 ();
 sg13g2_fill_2 FILLER_11_563 ();
 sg13g2_fill_2 FILLER_11_592 ();
 sg13g2_fill_2 FILLER_11_655 ();
 sg13g2_fill_2 FILLER_11_665 ();
 sg13g2_fill_2 FILLER_11_682 ();
 sg13g2_fill_1 FILLER_11_747 ();
 sg13g2_fill_2 FILLER_11_786 ();
 sg13g2_fill_2 FILLER_11_805 ();
 sg13g2_fill_2 FILLER_11_824 ();
 sg13g2_fill_1 FILLER_11_826 ();
 sg13g2_fill_2 FILLER_11_841 ();
 sg13g2_decap_8 FILLER_11_870 ();
 sg13g2_decap_8 FILLER_11_877 ();
 sg13g2_decap_8 FILLER_11_884 ();
 sg13g2_decap_8 FILLER_11_891 ();
 sg13g2_decap_8 FILLER_11_898 ();
 sg13g2_decap_8 FILLER_11_905 ();
 sg13g2_decap_8 FILLER_11_912 ();
 sg13g2_decap_8 FILLER_11_919 ();
 sg13g2_decap_8 FILLER_11_926 ();
 sg13g2_decap_8 FILLER_11_933 ();
 sg13g2_decap_8 FILLER_11_940 ();
 sg13g2_decap_8 FILLER_11_947 ();
 sg13g2_decap_8 FILLER_11_954 ();
 sg13g2_decap_8 FILLER_11_961 ();
 sg13g2_decap_8 FILLER_11_968 ();
 sg13g2_decap_8 FILLER_11_975 ();
 sg13g2_decap_8 FILLER_11_982 ();
 sg13g2_decap_8 FILLER_11_989 ();
 sg13g2_decap_8 FILLER_11_996 ();
 sg13g2_decap_8 FILLER_11_1003 ();
 sg13g2_decap_8 FILLER_11_1010 ();
 sg13g2_decap_8 FILLER_11_1017 ();
 sg13g2_decap_4 FILLER_11_1024 ();
 sg13g2_fill_1 FILLER_11_1028 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_282 ();
 sg13g2_fill_1 FILLER_12_297 ();
 sg13g2_fill_1 FILLER_12_315 ();
 sg13g2_fill_2 FILLER_12_330 ();
 sg13g2_fill_2 FILLER_12_341 ();
 sg13g2_fill_1 FILLER_12_343 ();
 sg13g2_fill_1 FILLER_12_371 ();
 sg13g2_fill_2 FILLER_12_395 ();
 sg13g2_fill_1 FILLER_12_434 ();
 sg13g2_fill_2 FILLER_12_461 ();
 sg13g2_fill_2 FILLER_12_467 ();
 sg13g2_fill_1 FILLER_12_469 ();
 sg13g2_fill_1 FILLER_12_510 ();
 sg13g2_fill_2 FILLER_12_548 ();
 sg13g2_fill_1 FILLER_12_550 ();
 sg13g2_fill_1 FILLER_12_586 ();
 sg13g2_fill_1 FILLER_12_636 ();
 sg13g2_fill_2 FILLER_12_666 ();
 sg13g2_fill_1 FILLER_12_668 ();
 sg13g2_fill_2 FILLER_12_774 ();
 sg13g2_fill_2 FILLER_12_802 ();
 sg13g2_fill_2 FILLER_12_824 ();
 sg13g2_decap_8 FILLER_12_865 ();
 sg13g2_decap_8 FILLER_12_872 ();
 sg13g2_decap_8 FILLER_12_879 ();
 sg13g2_decap_8 FILLER_12_886 ();
 sg13g2_decap_8 FILLER_12_893 ();
 sg13g2_decap_8 FILLER_12_900 ();
 sg13g2_decap_8 FILLER_12_907 ();
 sg13g2_decap_8 FILLER_12_914 ();
 sg13g2_decap_8 FILLER_12_921 ();
 sg13g2_decap_8 FILLER_12_928 ();
 sg13g2_decap_8 FILLER_12_935 ();
 sg13g2_decap_8 FILLER_12_942 ();
 sg13g2_decap_8 FILLER_12_949 ();
 sg13g2_decap_8 FILLER_12_956 ();
 sg13g2_decap_8 FILLER_12_963 ();
 sg13g2_decap_8 FILLER_12_970 ();
 sg13g2_decap_8 FILLER_12_977 ();
 sg13g2_decap_8 FILLER_12_984 ();
 sg13g2_decap_8 FILLER_12_991 ();
 sg13g2_decap_8 FILLER_12_998 ();
 sg13g2_decap_8 FILLER_12_1005 ();
 sg13g2_decap_8 FILLER_12_1012 ();
 sg13g2_decap_8 FILLER_12_1019 ();
 sg13g2_fill_2 FILLER_12_1026 ();
 sg13g2_fill_1 FILLER_12_1028 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_38 ();
 sg13g2_fill_1 FILLER_13_57 ();
 sg13g2_fill_1 FILLER_13_88 ();
 sg13g2_fill_2 FILLER_13_98 ();
 sg13g2_fill_2 FILLER_13_147 ();
 sg13g2_fill_1 FILLER_13_149 ();
 sg13g2_fill_2 FILLER_13_159 ();
 sg13g2_fill_1 FILLER_13_161 ();
 sg13g2_fill_2 FILLER_13_194 ();
 sg13g2_fill_2 FILLER_13_272 ();
 sg13g2_fill_2 FILLER_13_297 ();
 sg13g2_fill_1 FILLER_13_376 ();
 sg13g2_fill_2 FILLER_13_390 ();
 sg13g2_fill_2 FILLER_13_430 ();
 sg13g2_fill_1 FILLER_13_432 ();
 sg13g2_fill_2 FILLER_13_445 ();
 sg13g2_fill_1 FILLER_13_475 ();
 sg13g2_fill_2 FILLER_13_513 ();
 sg13g2_fill_1 FILLER_13_544 ();
 sg13g2_fill_1 FILLER_13_591 ();
 sg13g2_fill_2 FILLER_13_616 ();
 sg13g2_fill_2 FILLER_13_702 ();
 sg13g2_fill_1 FILLER_13_704 ();
 sg13g2_fill_2 FILLER_13_719 ();
 sg13g2_fill_1 FILLER_13_721 ();
 sg13g2_fill_1 FILLER_13_758 ();
 sg13g2_fill_1 FILLER_13_781 ();
 sg13g2_fill_1 FILLER_13_808 ();
 sg13g2_fill_1 FILLER_13_814 ();
 sg13g2_fill_1 FILLER_13_833 ();
 sg13g2_fill_2 FILLER_13_851 ();
 sg13g2_fill_1 FILLER_13_853 ();
 sg13g2_decap_8 FILLER_13_881 ();
 sg13g2_decap_8 FILLER_13_888 ();
 sg13g2_decap_8 FILLER_13_895 ();
 sg13g2_decap_8 FILLER_13_902 ();
 sg13g2_decap_8 FILLER_13_909 ();
 sg13g2_decap_8 FILLER_13_916 ();
 sg13g2_decap_8 FILLER_13_923 ();
 sg13g2_decap_8 FILLER_13_930 ();
 sg13g2_decap_8 FILLER_13_937 ();
 sg13g2_decap_8 FILLER_13_944 ();
 sg13g2_decap_8 FILLER_13_951 ();
 sg13g2_decap_8 FILLER_13_958 ();
 sg13g2_decap_8 FILLER_13_965 ();
 sg13g2_decap_8 FILLER_13_972 ();
 sg13g2_decap_8 FILLER_13_979 ();
 sg13g2_decap_8 FILLER_13_986 ();
 sg13g2_decap_8 FILLER_13_993 ();
 sg13g2_decap_8 FILLER_13_1000 ();
 sg13g2_decap_8 FILLER_13_1007 ();
 sg13g2_decap_8 FILLER_13_1014 ();
 sg13g2_decap_8 FILLER_13_1021 ();
 sg13g2_fill_1 FILLER_13_1028 ();
 sg13g2_fill_1 FILLER_14_118 ();
 sg13g2_fill_2 FILLER_14_142 ();
 sg13g2_fill_1 FILLER_14_144 ();
 sg13g2_fill_2 FILLER_14_159 ();
 sg13g2_fill_1 FILLER_14_187 ();
 sg13g2_fill_2 FILLER_14_290 ();
 sg13g2_fill_2 FILLER_14_418 ();
 sg13g2_fill_2 FILLER_14_437 ();
 sg13g2_fill_2 FILLER_14_448 ();
 sg13g2_fill_2 FILLER_14_526 ();
 sg13g2_decap_4 FILLER_14_582 ();
 sg13g2_fill_1 FILLER_14_603 ();
 sg13g2_fill_2 FILLER_14_637 ();
 sg13g2_fill_1 FILLER_14_639 ();
 sg13g2_fill_2 FILLER_14_690 ();
 sg13g2_fill_1 FILLER_14_692 ();
 sg13g2_fill_1 FILLER_14_734 ();
 sg13g2_fill_2 FILLER_14_758 ();
 sg13g2_fill_2 FILLER_14_779 ();
 sg13g2_fill_1 FILLER_14_790 ();
 sg13g2_fill_1 FILLER_14_850 ();
 sg13g2_decap_8 FILLER_14_878 ();
 sg13g2_decap_8 FILLER_14_885 ();
 sg13g2_decap_8 FILLER_14_892 ();
 sg13g2_decap_8 FILLER_14_899 ();
 sg13g2_decap_8 FILLER_14_906 ();
 sg13g2_decap_8 FILLER_14_913 ();
 sg13g2_decap_8 FILLER_14_920 ();
 sg13g2_decap_8 FILLER_14_927 ();
 sg13g2_decap_8 FILLER_14_934 ();
 sg13g2_decap_8 FILLER_14_941 ();
 sg13g2_decap_8 FILLER_14_948 ();
 sg13g2_decap_8 FILLER_14_955 ();
 sg13g2_decap_8 FILLER_14_962 ();
 sg13g2_decap_8 FILLER_14_969 ();
 sg13g2_decap_8 FILLER_14_976 ();
 sg13g2_decap_8 FILLER_14_983 ();
 sg13g2_decap_8 FILLER_14_990 ();
 sg13g2_decap_8 FILLER_14_997 ();
 sg13g2_decap_8 FILLER_14_1004 ();
 sg13g2_decap_8 FILLER_14_1011 ();
 sg13g2_decap_8 FILLER_14_1018 ();
 sg13g2_decap_4 FILLER_14_1025 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_193 ();
 sg13g2_fill_2 FILLER_15_223 ();
 sg13g2_fill_1 FILLER_15_225 ();
 sg13g2_fill_1 FILLER_15_259 ();
 sg13g2_fill_1 FILLER_15_404 ();
 sg13g2_fill_2 FILLER_15_439 ();
 sg13g2_fill_1 FILLER_15_441 ();
 sg13g2_fill_1 FILLER_15_533 ();
 sg13g2_fill_2 FILLER_15_539 ();
 sg13g2_decap_4 FILLER_15_577 ();
 sg13g2_fill_2 FILLER_15_627 ();
 sg13g2_fill_1 FILLER_15_629 ();
 sg13g2_fill_1 FILLER_15_714 ();
 sg13g2_fill_2 FILLER_15_756 ();
 sg13g2_fill_1 FILLER_15_787 ();
 sg13g2_fill_2 FILLER_15_798 ();
 sg13g2_fill_1 FILLER_15_845 ();
 sg13g2_decap_8 FILLER_15_885 ();
 sg13g2_decap_8 FILLER_15_892 ();
 sg13g2_decap_8 FILLER_15_899 ();
 sg13g2_decap_8 FILLER_15_906 ();
 sg13g2_decap_8 FILLER_15_913 ();
 sg13g2_decap_8 FILLER_15_920 ();
 sg13g2_decap_8 FILLER_15_927 ();
 sg13g2_decap_8 FILLER_15_934 ();
 sg13g2_decap_8 FILLER_15_941 ();
 sg13g2_decap_8 FILLER_15_948 ();
 sg13g2_decap_8 FILLER_15_955 ();
 sg13g2_decap_8 FILLER_15_962 ();
 sg13g2_decap_8 FILLER_15_969 ();
 sg13g2_decap_8 FILLER_15_976 ();
 sg13g2_decap_8 FILLER_15_983 ();
 sg13g2_decap_8 FILLER_15_990 ();
 sg13g2_decap_8 FILLER_15_997 ();
 sg13g2_decap_8 FILLER_15_1004 ();
 sg13g2_decap_8 FILLER_15_1011 ();
 sg13g2_decap_8 FILLER_15_1018 ();
 sg13g2_decap_4 FILLER_15_1025 ();
 sg13g2_fill_1 FILLER_16_32 ();
 sg13g2_fill_1 FILLER_16_74 ();
 sg13g2_fill_1 FILLER_16_84 ();
 sg13g2_fill_2 FILLER_16_148 ();
 sg13g2_fill_1 FILLER_16_194 ();
 sg13g2_fill_2 FILLER_16_272 ();
 sg13g2_fill_2 FILLER_16_353 ();
 sg13g2_fill_1 FILLER_16_405 ();
 sg13g2_fill_1 FILLER_16_415 ();
 sg13g2_fill_2 FILLER_16_430 ();
 sg13g2_fill_1 FILLER_16_522 ();
 sg13g2_fill_2 FILLER_16_536 ();
 sg13g2_fill_1 FILLER_16_547 ();
 sg13g2_decap_4 FILLER_16_576 ();
 sg13g2_fill_1 FILLER_16_580 ();
 sg13g2_fill_2 FILLER_16_683 ();
 sg13g2_fill_1 FILLER_16_744 ();
 sg13g2_fill_1 FILLER_16_750 ();
 sg13g2_fill_1 FILLER_16_803 ();
 sg13g2_fill_1 FILLER_16_870 ();
 sg13g2_fill_1 FILLER_16_880 ();
 sg13g2_decap_8 FILLER_16_886 ();
 sg13g2_decap_8 FILLER_16_893 ();
 sg13g2_decap_8 FILLER_16_900 ();
 sg13g2_decap_8 FILLER_16_907 ();
 sg13g2_decap_8 FILLER_16_914 ();
 sg13g2_decap_8 FILLER_16_921 ();
 sg13g2_decap_8 FILLER_16_928 ();
 sg13g2_decap_8 FILLER_16_935 ();
 sg13g2_decap_8 FILLER_16_942 ();
 sg13g2_decap_8 FILLER_16_949 ();
 sg13g2_decap_8 FILLER_16_956 ();
 sg13g2_decap_8 FILLER_16_963 ();
 sg13g2_decap_8 FILLER_16_970 ();
 sg13g2_decap_8 FILLER_16_977 ();
 sg13g2_decap_8 FILLER_16_984 ();
 sg13g2_decap_8 FILLER_16_991 ();
 sg13g2_decap_8 FILLER_16_998 ();
 sg13g2_decap_8 FILLER_16_1005 ();
 sg13g2_decap_8 FILLER_16_1012 ();
 sg13g2_decap_8 FILLER_16_1019 ();
 sg13g2_fill_2 FILLER_16_1026 ();
 sg13g2_fill_1 FILLER_16_1028 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_132 ();
 sg13g2_fill_2 FILLER_17_146 ();
 sg13g2_fill_1 FILLER_17_222 ();
 sg13g2_fill_2 FILLER_17_252 ();
 sg13g2_fill_1 FILLER_17_277 ();
 sg13g2_fill_1 FILLER_17_287 ();
 sg13g2_fill_2 FILLER_17_313 ();
 sg13g2_fill_2 FILLER_17_322 ();
 sg13g2_fill_1 FILLER_17_324 ();
 sg13g2_fill_1 FILLER_17_343 ();
 sg13g2_fill_1 FILLER_17_372 ();
 sg13g2_fill_2 FILLER_17_382 ();
 sg13g2_fill_1 FILLER_17_439 ();
 sg13g2_fill_1 FILLER_17_517 ();
 sg13g2_decap_4 FILLER_17_585 ();
 sg13g2_fill_1 FILLER_17_589 ();
 sg13g2_fill_1 FILLER_17_630 ();
 sg13g2_fill_2 FILLER_17_639 ();
 sg13g2_fill_1 FILLER_17_641 ();
 sg13g2_fill_1 FILLER_17_679 ();
 sg13g2_fill_2 FILLER_17_694 ();
 sg13g2_fill_1 FILLER_17_750 ();
 sg13g2_fill_1 FILLER_17_756 ();
 sg13g2_fill_1 FILLER_17_812 ();
 sg13g2_fill_2 FILLER_17_835 ();
 sg13g2_fill_2 FILLER_17_870 ();
 sg13g2_decap_8 FILLER_17_899 ();
 sg13g2_decap_8 FILLER_17_906 ();
 sg13g2_decap_8 FILLER_17_913 ();
 sg13g2_decap_8 FILLER_17_920 ();
 sg13g2_decap_8 FILLER_17_927 ();
 sg13g2_decap_8 FILLER_17_934 ();
 sg13g2_decap_8 FILLER_17_941 ();
 sg13g2_decap_8 FILLER_17_948 ();
 sg13g2_decap_8 FILLER_17_955 ();
 sg13g2_decap_8 FILLER_17_962 ();
 sg13g2_decap_8 FILLER_17_969 ();
 sg13g2_decap_8 FILLER_17_976 ();
 sg13g2_decap_8 FILLER_17_983 ();
 sg13g2_decap_8 FILLER_17_990 ();
 sg13g2_decap_8 FILLER_17_997 ();
 sg13g2_decap_8 FILLER_17_1004 ();
 sg13g2_decap_8 FILLER_17_1011 ();
 sg13g2_decap_8 FILLER_17_1018 ();
 sg13g2_decap_4 FILLER_17_1025 ();
 sg13g2_fill_2 FILLER_18_41 ();
 sg13g2_fill_1 FILLER_18_43 ();
 sg13g2_fill_1 FILLER_18_53 ();
 sg13g2_fill_2 FILLER_18_93 ();
 sg13g2_fill_1 FILLER_18_95 ();
 sg13g2_fill_2 FILLER_18_118 ();
 sg13g2_fill_1 FILLER_18_156 ();
 sg13g2_fill_2 FILLER_18_171 ();
 sg13g2_fill_2 FILLER_18_186 ();
 sg13g2_fill_1 FILLER_18_220 ();
 sg13g2_fill_1 FILLER_18_306 ();
 sg13g2_fill_2 FILLER_18_397 ();
 sg13g2_fill_1 FILLER_18_399 ();
 sg13g2_fill_1 FILLER_18_414 ();
 sg13g2_fill_2 FILLER_18_440 ();
 sg13g2_fill_1 FILLER_18_442 ();
 sg13g2_fill_2 FILLER_18_456 ();
 sg13g2_fill_1 FILLER_18_458 ();
 sg13g2_fill_2 FILLER_18_487 ();
 sg13g2_fill_2 FILLER_18_518 ();
 sg13g2_fill_1 FILLER_18_537 ();
 sg13g2_fill_1 FILLER_18_552 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_4 FILLER_18_588 ();
 sg13g2_fill_2 FILLER_18_671 ();
 sg13g2_fill_1 FILLER_18_683 ();
 sg13g2_fill_2 FILLER_18_714 ();
 sg13g2_fill_1 FILLER_18_729 ();
 sg13g2_fill_2 FILLER_18_760 ();
 sg13g2_fill_1 FILLER_18_822 ();
 sg13g2_fill_2 FILLER_18_851 ();
 sg13g2_fill_1 FILLER_18_872 ();
 sg13g2_decap_8 FILLER_18_905 ();
 sg13g2_decap_8 FILLER_18_912 ();
 sg13g2_decap_8 FILLER_18_919 ();
 sg13g2_decap_8 FILLER_18_926 ();
 sg13g2_decap_8 FILLER_18_933 ();
 sg13g2_decap_8 FILLER_18_940 ();
 sg13g2_decap_8 FILLER_18_947 ();
 sg13g2_decap_8 FILLER_18_954 ();
 sg13g2_decap_8 FILLER_18_961 ();
 sg13g2_decap_8 FILLER_18_968 ();
 sg13g2_decap_8 FILLER_18_975 ();
 sg13g2_decap_8 FILLER_18_982 ();
 sg13g2_decap_8 FILLER_18_989 ();
 sg13g2_decap_8 FILLER_18_996 ();
 sg13g2_decap_8 FILLER_18_1003 ();
 sg13g2_decap_8 FILLER_18_1010 ();
 sg13g2_decap_8 FILLER_18_1017 ();
 sg13g2_decap_4 FILLER_18_1024 ();
 sg13g2_fill_1 FILLER_18_1028 ();
 sg13g2_fill_1 FILLER_19_77 ();
 sg13g2_fill_2 FILLER_19_105 ();
 sg13g2_fill_1 FILLER_19_107 ();
 sg13g2_fill_1 FILLER_19_125 ();
 sg13g2_fill_1 FILLER_19_145 ();
 sg13g2_fill_2 FILLER_19_154 ();
 sg13g2_fill_1 FILLER_19_156 ();
 sg13g2_fill_1 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_217 ();
 sg13g2_fill_1 FILLER_19_278 ();
 sg13g2_fill_1 FILLER_19_298 ();
 sg13g2_fill_1 FILLER_19_319 ();
 sg13g2_fill_2 FILLER_19_348 ();
 sg13g2_fill_2 FILLER_19_422 ();
 sg13g2_fill_1 FILLER_19_424 ();
 sg13g2_fill_1 FILLER_19_447 ();
 sg13g2_fill_1 FILLER_19_494 ();
 sg13g2_fill_1 FILLER_19_508 ();
 sg13g2_fill_1 FILLER_19_683 ();
 sg13g2_fill_1 FILLER_19_780 ();
 sg13g2_fill_1 FILLER_19_804 ();
 sg13g2_fill_2 FILLER_19_837 ();
 sg13g2_fill_2 FILLER_19_849 ();
 sg13g2_decap_8 FILLER_19_912 ();
 sg13g2_decap_8 FILLER_19_919 ();
 sg13g2_decap_8 FILLER_19_926 ();
 sg13g2_decap_8 FILLER_19_933 ();
 sg13g2_decap_8 FILLER_19_940 ();
 sg13g2_decap_8 FILLER_19_947 ();
 sg13g2_decap_8 FILLER_19_954 ();
 sg13g2_decap_8 FILLER_19_961 ();
 sg13g2_decap_8 FILLER_19_968 ();
 sg13g2_decap_8 FILLER_19_975 ();
 sg13g2_decap_8 FILLER_19_982 ();
 sg13g2_decap_8 FILLER_19_989 ();
 sg13g2_decap_8 FILLER_19_996 ();
 sg13g2_decap_8 FILLER_19_1003 ();
 sg13g2_decap_8 FILLER_19_1010 ();
 sg13g2_decap_8 FILLER_19_1017 ();
 sg13g2_decap_4 FILLER_19_1024 ();
 sg13g2_fill_1 FILLER_19_1028 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_fill_2 FILLER_20_79 ();
 sg13g2_fill_1 FILLER_20_81 ();
 sg13g2_fill_2 FILLER_20_118 ();
 sg13g2_fill_1 FILLER_20_142 ();
 sg13g2_fill_1 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_343 ();
 sg13g2_fill_1 FILLER_20_345 ();
 sg13g2_fill_2 FILLER_20_374 ();
 sg13g2_fill_1 FILLER_20_376 ();
 sg13g2_fill_2 FILLER_20_396 ();
 sg13g2_fill_2 FILLER_20_408 ();
 sg13g2_fill_2 FILLER_20_423 ();
 sg13g2_fill_1 FILLER_20_425 ();
 sg13g2_fill_1 FILLER_20_492 ();
 sg13g2_fill_2 FILLER_20_551 ();
 sg13g2_fill_1 FILLER_20_553 ();
 sg13g2_fill_2 FILLER_20_639 ();
 sg13g2_fill_1 FILLER_20_641 ();
 sg13g2_fill_2 FILLER_20_829 ();
 sg13g2_decap_8 FILLER_20_919 ();
 sg13g2_decap_8 FILLER_20_926 ();
 sg13g2_decap_8 FILLER_20_933 ();
 sg13g2_decap_8 FILLER_20_940 ();
 sg13g2_decap_8 FILLER_20_947 ();
 sg13g2_decap_8 FILLER_20_954 ();
 sg13g2_decap_8 FILLER_20_961 ();
 sg13g2_decap_8 FILLER_20_968 ();
 sg13g2_decap_8 FILLER_20_975 ();
 sg13g2_decap_8 FILLER_20_982 ();
 sg13g2_decap_8 FILLER_20_989 ();
 sg13g2_decap_8 FILLER_20_996 ();
 sg13g2_decap_8 FILLER_20_1003 ();
 sg13g2_decap_8 FILLER_20_1010 ();
 sg13g2_decap_8 FILLER_20_1017 ();
 sg13g2_decap_4 FILLER_20_1024 ();
 sg13g2_fill_1 FILLER_20_1028 ();
 sg13g2_fill_2 FILLER_21_60 ();
 sg13g2_fill_2 FILLER_21_76 ();
 sg13g2_fill_1 FILLER_21_106 ();
 sg13g2_fill_1 FILLER_21_143 ();
 sg13g2_fill_1 FILLER_21_160 ();
 sg13g2_fill_1 FILLER_21_178 ();
 sg13g2_fill_1 FILLER_21_314 ();
 sg13g2_fill_1 FILLER_21_324 ();
 sg13g2_fill_2 FILLER_21_347 ();
 sg13g2_fill_1 FILLER_21_349 ();
 sg13g2_fill_2 FILLER_21_385 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_2 FILLER_21_451 ();
 sg13g2_fill_2 FILLER_21_477 ();
 sg13g2_fill_1 FILLER_21_483 ();
 sg13g2_fill_1 FILLER_21_511 ();
 sg13g2_fill_1 FILLER_21_525 ();
 sg13g2_fill_2 FILLER_21_570 ();
 sg13g2_fill_1 FILLER_21_580 ();
 sg13g2_fill_2 FILLER_21_742 ();
 sg13g2_fill_1 FILLER_21_784 ();
 sg13g2_fill_1 FILLER_21_798 ();
 sg13g2_fill_1 FILLER_21_812 ();
 sg13g2_fill_1 FILLER_21_858 ();
 sg13g2_fill_2 FILLER_21_910 ();
 sg13g2_decap_8 FILLER_21_926 ();
 sg13g2_decap_8 FILLER_21_933 ();
 sg13g2_decap_8 FILLER_21_940 ();
 sg13g2_decap_8 FILLER_21_947 ();
 sg13g2_decap_8 FILLER_21_954 ();
 sg13g2_decap_8 FILLER_21_961 ();
 sg13g2_decap_8 FILLER_21_968 ();
 sg13g2_decap_8 FILLER_21_975 ();
 sg13g2_decap_8 FILLER_21_982 ();
 sg13g2_decap_8 FILLER_21_989 ();
 sg13g2_decap_8 FILLER_21_996 ();
 sg13g2_decap_8 FILLER_21_1003 ();
 sg13g2_decap_8 FILLER_21_1010 ();
 sg13g2_decap_8 FILLER_21_1017 ();
 sg13g2_decap_4 FILLER_21_1024 ();
 sg13g2_fill_1 FILLER_21_1028 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_fill_1 FILLER_22_70 ();
 sg13g2_fill_1 FILLER_22_166 ();
 sg13g2_fill_1 FILLER_22_197 ();
 sg13g2_fill_2 FILLER_22_262 ();
 sg13g2_fill_2 FILLER_22_334 ();
 sg13g2_fill_2 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_510 ();
 sg13g2_fill_1 FILLER_22_529 ();
 sg13g2_fill_1 FILLER_22_539 ();
 sg13g2_decap_4 FILLER_22_608 ();
 sg13g2_fill_2 FILLER_22_627 ();
 sg13g2_fill_2 FILLER_22_666 ();
 sg13g2_fill_1 FILLER_22_668 ();
 sg13g2_fill_1 FILLER_22_679 ();
 sg13g2_fill_2 FILLER_22_780 ();
 sg13g2_fill_1 FILLER_22_827 ();
 sg13g2_fill_2 FILLER_22_850 ();
 sg13g2_fill_2 FILLER_22_884 ();
 sg13g2_decap_8 FILLER_22_923 ();
 sg13g2_decap_8 FILLER_22_930 ();
 sg13g2_decap_8 FILLER_22_937 ();
 sg13g2_decap_8 FILLER_22_944 ();
 sg13g2_decap_8 FILLER_22_951 ();
 sg13g2_decap_8 FILLER_22_958 ();
 sg13g2_decap_8 FILLER_22_965 ();
 sg13g2_decap_8 FILLER_22_972 ();
 sg13g2_decap_8 FILLER_22_979 ();
 sg13g2_decap_8 FILLER_22_986 ();
 sg13g2_decap_8 FILLER_22_993 ();
 sg13g2_decap_8 FILLER_22_1000 ();
 sg13g2_decap_8 FILLER_22_1007 ();
 sg13g2_decap_8 FILLER_22_1014 ();
 sg13g2_decap_8 FILLER_22_1021 ();
 sg13g2_fill_1 FILLER_22_1028 ();
 sg13g2_fill_2 FILLER_23_108 ();
 sg13g2_fill_1 FILLER_23_140 ();
 sg13g2_fill_2 FILLER_23_148 ();
 sg13g2_fill_1 FILLER_23_166 ();
 sg13g2_fill_1 FILLER_23_237 ();
 sg13g2_fill_1 FILLER_23_251 ();
 sg13g2_fill_2 FILLER_23_261 ();
 sg13g2_fill_1 FILLER_23_277 ();
 sg13g2_fill_2 FILLER_23_317 ();
 sg13g2_fill_1 FILLER_23_319 ();
 sg13g2_fill_2 FILLER_23_343 ();
 sg13g2_fill_1 FILLER_23_381 ();
 sg13g2_fill_2 FILLER_23_451 ();
 sg13g2_fill_1 FILLER_23_481 ();
 sg13g2_fill_2 FILLER_23_527 ();
 sg13g2_fill_1 FILLER_23_538 ();
 sg13g2_fill_1 FILLER_23_548 ();
 sg13g2_fill_1 FILLER_23_562 ();
 sg13g2_fill_2 FILLER_23_661 ();
 sg13g2_fill_1 FILLER_23_676 ();
 sg13g2_fill_2 FILLER_23_705 ();
 sg13g2_fill_1 FILLER_23_707 ();
 sg13g2_fill_2 FILLER_23_763 ();
 sg13g2_fill_1 FILLER_23_794 ();
 sg13g2_fill_1 FILLER_23_800 ();
 sg13g2_fill_2 FILLER_23_858 ();
 sg13g2_fill_2 FILLER_23_878 ();
 sg13g2_decap_8 FILLER_23_922 ();
 sg13g2_decap_8 FILLER_23_929 ();
 sg13g2_decap_8 FILLER_23_936 ();
 sg13g2_decap_8 FILLER_23_943 ();
 sg13g2_decap_8 FILLER_23_950 ();
 sg13g2_decap_8 FILLER_23_957 ();
 sg13g2_decap_8 FILLER_23_964 ();
 sg13g2_decap_8 FILLER_23_971 ();
 sg13g2_decap_8 FILLER_23_978 ();
 sg13g2_decap_8 FILLER_23_985 ();
 sg13g2_decap_8 FILLER_23_992 ();
 sg13g2_decap_8 FILLER_23_999 ();
 sg13g2_decap_8 FILLER_23_1006 ();
 sg13g2_decap_8 FILLER_23_1013 ();
 sg13g2_decap_8 FILLER_23_1020 ();
 sg13g2_fill_2 FILLER_23_1027 ();
 sg13g2_fill_2 FILLER_24_40 ();
 sg13g2_fill_1 FILLER_24_42 ();
 sg13g2_fill_1 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_73 ();
 sg13g2_fill_1 FILLER_24_129 ();
 sg13g2_fill_1 FILLER_24_165 ();
 sg13g2_fill_2 FILLER_24_200 ();
 sg13g2_fill_1 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_251 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_fill_1 FILLER_24_285 ();
 sg13g2_fill_2 FILLER_24_343 ();
 sg13g2_fill_1 FILLER_24_345 ();
 sg13g2_fill_2 FILLER_24_381 ();
 sg13g2_fill_1 FILLER_24_383 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_fill_2 FILLER_24_444 ();
 sg13g2_fill_1 FILLER_24_489 ();
 sg13g2_fill_1 FILLER_24_512 ();
 sg13g2_fill_1 FILLER_24_550 ();
 sg13g2_fill_2 FILLER_24_640 ();
 sg13g2_fill_2 FILLER_24_696 ();
 sg13g2_fill_1 FILLER_24_698 ();
 sg13g2_fill_1 FILLER_24_747 ();
 sg13g2_fill_1 FILLER_24_787 ();
 sg13g2_fill_2 FILLER_24_819 ();
 sg13g2_fill_2 FILLER_24_829 ();
 sg13g2_fill_1 FILLER_24_868 ();
 sg13g2_fill_1 FILLER_24_884 ();
 sg13g2_fill_2 FILLER_24_890 ();
 sg13g2_fill_1 FILLER_24_933 ();
 sg13g2_decap_8 FILLER_24_946 ();
 sg13g2_decap_8 FILLER_24_953 ();
 sg13g2_decap_8 FILLER_24_960 ();
 sg13g2_decap_8 FILLER_24_967 ();
 sg13g2_decap_8 FILLER_24_974 ();
 sg13g2_decap_8 FILLER_24_981 ();
 sg13g2_decap_8 FILLER_24_988 ();
 sg13g2_decap_8 FILLER_24_995 ();
 sg13g2_decap_8 FILLER_24_1002 ();
 sg13g2_decap_8 FILLER_24_1009 ();
 sg13g2_decap_8 FILLER_24_1016 ();
 sg13g2_decap_4 FILLER_24_1023 ();
 sg13g2_fill_2 FILLER_24_1027 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_40 ();
 sg13g2_fill_2 FILLER_25_103 ();
 sg13g2_fill_1 FILLER_25_109 ();
 sg13g2_fill_1 FILLER_25_129 ();
 sg13g2_fill_1 FILLER_25_138 ();
 sg13g2_fill_2 FILLER_25_187 ();
 sg13g2_fill_2 FILLER_25_194 ();
 sg13g2_fill_1 FILLER_25_204 ();
 sg13g2_fill_2 FILLER_25_215 ();
 sg13g2_fill_2 FILLER_25_286 ();
 sg13g2_fill_2 FILLER_25_316 ();
 sg13g2_fill_2 FILLER_25_342 ();
 sg13g2_fill_2 FILLER_25_371 ();
 sg13g2_fill_1 FILLER_25_415 ();
 sg13g2_fill_2 FILLER_25_518 ();
 sg13g2_fill_2 FILLER_25_621 ();
 sg13g2_fill_1 FILLER_25_654 ();
 sg13g2_fill_2 FILLER_25_675 ();
 sg13g2_fill_1 FILLER_25_677 ();
 sg13g2_fill_1 FILLER_25_736 ();
 sg13g2_fill_2 FILLER_25_741 ();
 sg13g2_fill_1 FILLER_25_773 ();
 sg13g2_fill_1 FILLER_25_808 ();
 sg13g2_fill_2 FILLER_25_853 ();
 sg13g2_fill_1 FILLER_25_945 ();
 sg13g2_decap_8 FILLER_25_954 ();
 sg13g2_decap_8 FILLER_25_961 ();
 sg13g2_decap_8 FILLER_25_968 ();
 sg13g2_decap_8 FILLER_25_975 ();
 sg13g2_decap_8 FILLER_25_982 ();
 sg13g2_decap_8 FILLER_25_989 ();
 sg13g2_decap_8 FILLER_25_996 ();
 sg13g2_decap_8 FILLER_25_1003 ();
 sg13g2_decap_8 FILLER_25_1010 ();
 sg13g2_decap_8 FILLER_25_1017 ();
 sg13g2_decap_4 FILLER_25_1024 ();
 sg13g2_fill_1 FILLER_25_1028 ();
 sg13g2_fill_1 FILLER_26_12 ();
 sg13g2_fill_1 FILLER_26_52 ();
 sg13g2_fill_1 FILLER_26_61 ();
 sg13g2_fill_1 FILLER_26_107 ();
 sg13g2_fill_1 FILLER_26_125 ();
 sg13g2_fill_1 FILLER_26_139 ();
 sg13g2_fill_1 FILLER_26_145 ();
 sg13g2_fill_2 FILLER_26_162 ();
 sg13g2_fill_2 FILLER_26_172 ();
 sg13g2_fill_2 FILLER_26_187 ();
 sg13g2_fill_2 FILLER_26_222 ();
 sg13g2_fill_2 FILLER_26_256 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_fill_1 FILLER_26_313 ();
 sg13g2_fill_1 FILLER_26_322 ();
 sg13g2_fill_2 FILLER_26_339 ();
 sg13g2_fill_1 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_419 ();
 sg13g2_fill_1 FILLER_26_421 ();
 sg13g2_fill_2 FILLER_26_434 ();
 sg13g2_fill_1 FILLER_26_463 ();
 sg13g2_fill_2 FILLER_26_487 ();
 sg13g2_fill_2 FILLER_26_518 ();
 sg13g2_decap_8 FILLER_26_623 ();
 sg13g2_fill_2 FILLER_26_630 ();
 sg13g2_fill_1 FILLER_26_645 ();
 sg13g2_fill_1 FILLER_26_686 ();
 sg13g2_fill_2 FILLER_26_760 ();
 sg13g2_fill_1 FILLER_26_772 ();
 sg13g2_fill_2 FILLER_26_788 ();
 sg13g2_fill_2 FILLER_26_807 ();
 sg13g2_fill_2 FILLER_26_822 ();
 sg13g2_fill_1 FILLER_26_824 ();
 sg13g2_fill_1 FILLER_26_835 ();
 sg13g2_fill_1 FILLER_26_862 ();
 sg13g2_fill_1 FILLER_26_908 ();
 sg13g2_fill_1 FILLER_26_936 ();
 sg13g2_fill_1 FILLER_26_956 ();
 sg13g2_decap_8 FILLER_26_965 ();
 sg13g2_decap_8 FILLER_26_972 ();
 sg13g2_decap_8 FILLER_26_979 ();
 sg13g2_decap_8 FILLER_26_986 ();
 sg13g2_decap_8 FILLER_26_993 ();
 sg13g2_decap_8 FILLER_26_1000 ();
 sg13g2_decap_8 FILLER_26_1007 ();
 sg13g2_decap_8 FILLER_26_1014 ();
 sg13g2_decap_8 FILLER_26_1021 ();
 sg13g2_fill_1 FILLER_26_1028 ();
 sg13g2_fill_1 FILLER_27_4 ();
 sg13g2_fill_2 FILLER_27_37 ();
 sg13g2_fill_1 FILLER_27_39 ();
 sg13g2_fill_1 FILLER_27_69 ();
 sg13g2_fill_1 FILLER_27_125 ();
 sg13g2_fill_2 FILLER_27_162 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_219 ();
 sg13g2_fill_2 FILLER_27_236 ();
 sg13g2_fill_2 FILLER_27_362 ();
 sg13g2_fill_1 FILLER_27_364 ();
 sg13g2_fill_2 FILLER_27_414 ();
 sg13g2_fill_1 FILLER_27_416 ();
 sg13g2_fill_2 FILLER_27_448 ();
 sg13g2_fill_1 FILLER_27_503 ();
 sg13g2_fill_1 FILLER_27_514 ();
 sg13g2_fill_1 FILLER_27_550 ();
 sg13g2_fill_2 FILLER_27_625 ();
 sg13g2_fill_1 FILLER_27_627 ();
 sg13g2_fill_2 FILLER_27_659 ();
 sg13g2_fill_2 FILLER_27_764 ();
 sg13g2_fill_2 FILLER_27_782 ();
 sg13g2_fill_2 FILLER_27_806 ();
 sg13g2_fill_1 FILLER_27_825 ();
 sg13g2_fill_2 FILLER_27_844 ();
 sg13g2_fill_1 FILLER_27_846 ();
 sg13g2_fill_1 FILLER_27_856 ();
 sg13g2_decap_8 FILLER_27_974 ();
 sg13g2_decap_8 FILLER_27_981 ();
 sg13g2_decap_8 FILLER_27_988 ();
 sg13g2_decap_8 FILLER_27_995 ();
 sg13g2_decap_8 FILLER_27_1002 ();
 sg13g2_decap_8 FILLER_27_1009 ();
 sg13g2_decap_8 FILLER_27_1016 ();
 sg13g2_decap_4 FILLER_27_1023 ();
 sg13g2_fill_2 FILLER_27_1027 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_37 ();
 sg13g2_fill_1 FILLER_28_113 ();
 sg13g2_fill_2 FILLER_28_126 ();
 sg13g2_fill_1 FILLER_28_147 ();
 sg13g2_fill_1 FILLER_28_228 ();
 sg13g2_fill_2 FILLER_28_236 ();
 sg13g2_fill_2 FILLER_28_262 ();
 sg13g2_fill_2 FILLER_28_277 ();
 sg13g2_fill_2 FILLER_28_306 ();
 sg13g2_fill_1 FILLER_28_308 ();
 sg13g2_fill_2 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_444 ();
 sg13g2_fill_2 FILLER_28_478 ();
 sg13g2_fill_1 FILLER_28_548 ();
 sg13g2_fill_2 FILLER_28_589 ();
 sg13g2_fill_1 FILLER_28_591 ();
 sg13g2_fill_1 FILLER_28_637 ();
 sg13g2_fill_1 FILLER_28_661 ();
 sg13g2_fill_1 FILLER_28_690 ();
 sg13g2_fill_2 FILLER_28_774 ();
 sg13g2_fill_2 FILLER_28_780 ();
 sg13g2_fill_1 FILLER_28_808 ();
 sg13g2_fill_2 FILLER_28_846 ();
 sg13g2_fill_1 FILLER_28_848 ();
 sg13g2_fill_1 FILLER_28_928 ();
 sg13g2_decap_8 FILLER_28_985 ();
 sg13g2_decap_8 FILLER_28_992 ();
 sg13g2_decap_8 FILLER_28_999 ();
 sg13g2_decap_8 FILLER_28_1006 ();
 sg13g2_decap_8 FILLER_28_1013 ();
 sg13g2_decap_8 FILLER_28_1020 ();
 sg13g2_fill_2 FILLER_28_1027 ();
 sg13g2_fill_1 FILLER_29_8 ();
 sg13g2_fill_2 FILLER_29_36 ();
 sg13g2_fill_1 FILLER_29_38 ();
 sg13g2_fill_2 FILLER_29_65 ();
 sg13g2_fill_2 FILLER_29_107 ();
 sg13g2_fill_1 FILLER_29_126 ();
 sg13g2_fill_2 FILLER_29_192 ();
 sg13g2_fill_1 FILLER_29_194 ();
 sg13g2_fill_1 FILLER_29_207 ();
 sg13g2_fill_2 FILLER_29_232 ();
 sg13g2_fill_1 FILLER_29_256 ();
 sg13g2_fill_2 FILLER_29_294 ();
 sg13g2_fill_2 FILLER_29_340 ();
 sg13g2_fill_1 FILLER_29_342 ();
 sg13g2_fill_2 FILLER_29_361 ();
 sg13g2_fill_1 FILLER_29_447 ();
 sg13g2_fill_1 FILLER_29_470 ();
 sg13g2_fill_2 FILLER_29_481 ();
 sg13g2_fill_1 FILLER_29_510 ();
 sg13g2_decap_4 FILLER_29_527 ();
 sg13g2_fill_2 FILLER_29_531 ();
 sg13g2_fill_2 FILLER_29_571 ();
 sg13g2_fill_2 FILLER_29_587 ();
 sg13g2_fill_1 FILLER_29_589 ();
 sg13g2_fill_2 FILLER_29_644 ();
 sg13g2_fill_1 FILLER_29_646 ();
 sg13g2_fill_1 FILLER_29_703 ();
 sg13g2_fill_1 FILLER_29_786 ();
 sg13g2_fill_1 FILLER_29_808 ();
 sg13g2_fill_1 FILLER_29_822 ();
 sg13g2_fill_2 FILLER_29_827 ();
 sg13g2_fill_2 FILLER_29_897 ();
 sg13g2_fill_1 FILLER_29_899 ();
 sg13g2_decap_8 FILLER_29_997 ();
 sg13g2_decap_8 FILLER_29_1004 ();
 sg13g2_decap_8 FILLER_29_1011 ();
 sg13g2_decap_8 FILLER_29_1018 ();
 sg13g2_decap_4 FILLER_29_1025 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_fill_1 FILLER_30_50 ();
 sg13g2_fill_2 FILLER_30_59 ();
 sg13g2_fill_1 FILLER_30_61 ();
 sg13g2_fill_1 FILLER_30_69 ();
 sg13g2_fill_2 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_114 ();
 sg13g2_fill_1 FILLER_30_150 ();
 sg13g2_fill_1 FILLER_30_270 ();
 sg13g2_fill_2 FILLER_30_289 ();
 sg13g2_fill_2 FILLER_30_313 ();
 sg13g2_fill_1 FILLER_30_357 ();
 sg13g2_fill_2 FILLER_30_389 ();
 sg13g2_fill_1 FILLER_30_391 ();
 sg13g2_fill_2 FILLER_30_410 ();
 sg13g2_fill_1 FILLER_30_452 ();
 sg13g2_fill_1 FILLER_30_466 ();
 sg13g2_fill_2 FILLER_30_490 ();
 sg13g2_decap_8 FILLER_30_501 ();
 sg13g2_fill_1 FILLER_30_558 ();
 sg13g2_fill_2 FILLER_30_581 ();
 sg13g2_fill_1 FILLER_30_647 ();
 sg13g2_fill_2 FILLER_30_688 ();
 sg13g2_fill_2 FILLER_30_695 ();
 sg13g2_fill_1 FILLER_30_697 ();
 sg13g2_fill_2 FILLER_30_716 ();
 sg13g2_fill_1 FILLER_30_718 ();
 sg13g2_fill_2 FILLER_30_802 ();
 sg13g2_fill_1 FILLER_30_864 ();
 sg13g2_fill_1 FILLER_30_949 ();
 sg13g2_decap_8 FILLER_30_1006 ();
 sg13g2_decap_8 FILLER_30_1013 ();
 sg13g2_decap_8 FILLER_30_1020 ();
 sg13g2_fill_2 FILLER_30_1027 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_fill_1 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_27 ();
 sg13g2_fill_1 FILLER_31_96 ();
 sg13g2_fill_1 FILLER_31_110 ();
 sg13g2_fill_1 FILLER_31_161 ();
 sg13g2_fill_1 FILLER_31_204 ();
 sg13g2_fill_1 FILLER_31_258 ();
 sg13g2_fill_1 FILLER_31_332 ();
 sg13g2_fill_2 FILLER_31_351 ();
 sg13g2_fill_1 FILLER_31_353 ();
 sg13g2_fill_2 FILLER_31_421 ();
 sg13g2_fill_1 FILLER_31_423 ();
 sg13g2_fill_2 FILLER_31_437 ();
 sg13g2_fill_1 FILLER_31_439 ();
 sg13g2_fill_1 FILLER_31_481 ();
 sg13g2_decap_8 FILLER_31_498 ();
 sg13g2_fill_2 FILLER_31_571 ();
 sg13g2_fill_2 FILLER_31_597 ();
 sg13g2_fill_1 FILLER_31_599 ();
 sg13g2_fill_2 FILLER_31_628 ();
 sg13g2_fill_2 FILLER_31_674 ();
 sg13g2_fill_1 FILLER_31_676 ();
 sg13g2_fill_1 FILLER_31_691 ();
 sg13g2_fill_2 FILLER_31_762 ();
 sg13g2_fill_2 FILLER_31_769 ();
 sg13g2_fill_1 FILLER_31_789 ();
 sg13g2_fill_2 FILLER_31_798 ();
 sg13g2_fill_2 FILLER_31_895 ();
 sg13g2_fill_2 FILLER_31_936 ();
 sg13g2_fill_1 FILLER_31_991 ();
 sg13g2_decap_8 FILLER_31_1013 ();
 sg13g2_decap_8 FILLER_31_1020 ();
 sg13g2_fill_2 FILLER_31_1027 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_34 ();
 sg13g2_fill_1 FILLER_32_36 ();
 sg13g2_fill_2 FILLER_32_66 ();
 sg13g2_fill_1 FILLER_32_68 ();
 sg13g2_fill_2 FILLER_32_117 ();
 sg13g2_fill_1 FILLER_32_156 ();
 sg13g2_fill_2 FILLER_32_200 ();
 sg13g2_fill_1 FILLER_32_210 ();
 sg13g2_fill_1 FILLER_32_228 ();
 sg13g2_fill_1 FILLER_32_251 ();
 sg13g2_fill_1 FILLER_32_332 ();
 sg13g2_fill_2 FILLER_32_379 ();
 sg13g2_fill_2 FILLER_32_439 ();
 sg13g2_fill_1 FILLER_32_472 ();
 sg13g2_fill_2 FILLER_32_478 ();
 sg13g2_fill_1 FILLER_32_480 ();
 sg13g2_fill_2 FILLER_32_508 ();
 sg13g2_decap_4 FILLER_32_518 ();
 sg13g2_fill_2 FILLER_32_522 ();
 sg13g2_fill_1 FILLER_32_569 ();
 sg13g2_fill_2 FILLER_32_633 ();
 sg13g2_fill_1 FILLER_32_682 ();
 sg13g2_fill_2 FILLER_32_760 ();
 sg13g2_fill_2 FILLER_32_796 ();
 sg13g2_fill_1 FILLER_32_847 ();
 sg13g2_fill_2 FILLER_32_997 ();
 sg13g2_fill_2 FILLER_32_1026 ();
 sg13g2_fill_1 FILLER_32_1028 ();
 sg13g2_fill_1 FILLER_33_8 ();
 sg13g2_fill_2 FILLER_33_18 ();
 sg13g2_fill_1 FILLER_33_20 ();
 sg13g2_fill_1 FILLER_33_111 ();
 sg13g2_fill_2 FILLER_33_166 ();
 sg13g2_fill_1 FILLER_33_168 ();
 sg13g2_fill_2 FILLER_33_195 ();
 sg13g2_fill_1 FILLER_33_216 ();
 sg13g2_fill_2 FILLER_33_233 ();
 sg13g2_fill_1 FILLER_33_275 ();
 sg13g2_fill_2 FILLER_33_308 ();
 sg13g2_fill_2 FILLER_33_369 ();
 sg13g2_fill_1 FILLER_33_389 ();
 sg13g2_fill_1 FILLER_33_452 ();
 sg13g2_fill_2 FILLER_33_536 ();
 sg13g2_fill_1 FILLER_33_551 ();
 sg13g2_fill_1 FILLER_33_562 ();
 sg13g2_fill_2 FILLER_33_601 ();
 sg13g2_fill_1 FILLER_33_634 ();
 sg13g2_fill_2 FILLER_33_662 ();
 sg13g2_fill_2 FILLER_33_709 ();
 sg13g2_fill_2 FILLER_33_748 ();
 sg13g2_fill_1 FILLER_33_750 ();
 sg13g2_fill_1 FILLER_33_765 ();
 sg13g2_fill_1 FILLER_33_802 ();
 sg13g2_fill_1 FILLER_33_848 ();
 sg13g2_fill_1 FILLER_33_858 ();
 sg13g2_fill_1 FILLER_33_885 ();
 sg13g2_fill_1 FILLER_33_921 ();
 sg13g2_fill_1 FILLER_33_949 ();
 sg13g2_fill_1 FILLER_33_968 ();
 sg13g2_fill_1 FILLER_33_991 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_34 ();
 sg13g2_fill_2 FILLER_34_87 ();
 sg13g2_fill_1 FILLER_34_117 ();
 sg13g2_fill_1 FILLER_34_145 ();
 sg13g2_fill_1 FILLER_34_155 ();
 sg13g2_fill_2 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_192 ();
 sg13g2_fill_2 FILLER_34_217 ();
 sg13g2_fill_1 FILLER_34_219 ();
 sg13g2_fill_1 FILLER_34_237 ();
 sg13g2_fill_2 FILLER_34_271 ();
 sg13g2_fill_2 FILLER_34_321 ();
 sg13g2_fill_1 FILLER_34_323 ();
 sg13g2_fill_2 FILLER_34_382 ();
 sg13g2_fill_1 FILLER_34_456 ();
 sg13g2_fill_1 FILLER_34_474 ();
 sg13g2_fill_2 FILLER_34_498 ();
 sg13g2_decap_4 FILLER_34_528 ();
 sg13g2_fill_2 FILLER_34_581 ();
 sg13g2_fill_1 FILLER_34_596 ();
 sg13g2_fill_1 FILLER_34_629 ();
 sg13g2_fill_2 FILLER_34_744 ();
 sg13g2_fill_2 FILLER_34_766 ();
 sg13g2_fill_2 FILLER_34_827 ();
 sg13g2_fill_1 FILLER_34_829 ();
 sg13g2_fill_1 FILLER_34_843 ();
 sg13g2_fill_2 FILLER_34_970 ();
 sg13g2_fill_2 FILLER_34_985 ();
 sg13g2_fill_1 FILLER_34_987 ();
 sg13g2_fill_2 FILLER_34_993 ();
 sg13g2_fill_1 FILLER_34_995 ();
 sg13g2_fill_1 FILLER_35_8 ();
 sg13g2_fill_1 FILLER_35_26 ();
 sg13g2_fill_2 FILLER_35_51 ();
 sg13g2_fill_1 FILLER_35_53 ();
 sg13g2_fill_1 FILLER_35_86 ();
 sg13g2_fill_2 FILLER_35_114 ();
 sg13g2_fill_1 FILLER_35_116 ();
 sg13g2_fill_2 FILLER_35_232 ();
 sg13g2_fill_2 FILLER_35_269 ();
 sg13g2_fill_1 FILLER_35_271 ();
 sg13g2_fill_1 FILLER_35_303 ();
 sg13g2_fill_2 FILLER_35_313 ();
 sg13g2_fill_2 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_395 ();
 sg13g2_fill_2 FILLER_35_410 ();
 sg13g2_fill_2 FILLER_35_444 ();
 sg13g2_fill_1 FILLER_35_451 ();
 sg13g2_fill_1 FILLER_35_475 ();
 sg13g2_fill_2 FILLER_35_543 ();
 sg13g2_fill_1 FILLER_35_545 ();
 sg13g2_fill_2 FILLER_35_640 ();
 sg13g2_fill_1 FILLER_35_720 ();
 sg13g2_fill_1 FILLER_35_730 ();
 sg13g2_fill_2 FILLER_35_789 ();
 sg13g2_fill_1 FILLER_35_796 ();
 sg13g2_fill_2 FILLER_35_832 ();
 sg13g2_fill_2 FILLER_35_843 ();
 sg13g2_fill_2 FILLER_35_861 ();
 sg13g2_fill_2 FILLER_35_939 ();
 sg13g2_fill_2 FILLER_35_956 ();
 sg13g2_fill_2 FILLER_35_967 ();
 sg13g2_fill_2 FILLER_35_982 ();
 sg13g2_fill_1 FILLER_35_984 ();
 sg13g2_fill_2 FILLER_35_995 ();
 sg13g2_fill_2 FILLER_36_4 ();
 sg13g2_fill_2 FILLER_36_33 ();
 sg13g2_fill_1 FILLER_36_48 ();
 sg13g2_fill_1 FILLER_36_55 ();
 sg13g2_fill_1 FILLER_36_65 ();
 sg13g2_fill_1 FILLER_36_86 ();
 sg13g2_fill_1 FILLER_36_100 ();
 sg13g2_fill_1 FILLER_36_109 ();
 sg13g2_fill_2 FILLER_36_138 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_fill_2 FILLER_36_191 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_305 ();
 sg13g2_fill_1 FILLER_36_307 ();
 sg13g2_fill_1 FILLER_36_330 ();
 sg13g2_fill_1 FILLER_36_358 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_fill_2 FILLER_36_463 ();
 sg13g2_fill_2 FILLER_36_526 ();
 sg13g2_fill_2 FILLER_36_620 ();
 sg13g2_fill_1 FILLER_36_622 ();
 sg13g2_fill_1 FILLER_36_670 ();
 sg13g2_fill_1 FILLER_36_689 ();
 sg13g2_fill_1 FILLER_36_699 ();
 sg13g2_fill_2 FILLER_36_739 ();
 sg13g2_fill_2 FILLER_36_766 ();
 sg13g2_fill_2 FILLER_36_803 ();
 sg13g2_fill_2 FILLER_36_815 ();
 sg13g2_fill_1 FILLER_36_843 ();
 sg13g2_fill_2 FILLER_36_892 ();
 sg13g2_fill_1 FILLER_36_920 ();
 sg13g2_fill_2 FILLER_36_948 ();
 sg13g2_fill_1 FILLER_36_950 ();
 sg13g2_fill_2 FILLER_36_987 ();
 sg13g2_fill_1 FILLER_36_989 ();
 sg13g2_fill_1 FILLER_36_1017 ();
 sg13g2_fill_2 FILLER_36_1027 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_134 ();
 sg13g2_fill_2 FILLER_37_169 ();
 sg13g2_fill_1 FILLER_37_192 ();
 sg13g2_fill_2 FILLER_37_214 ();
 sg13g2_fill_1 FILLER_37_216 ();
 sg13g2_fill_1 FILLER_37_264 ();
 sg13g2_fill_2 FILLER_37_368 ();
 sg13g2_fill_1 FILLER_37_370 ();
 sg13g2_fill_2 FILLER_37_397 ();
 sg13g2_fill_1 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_422 ();
 sg13g2_fill_1 FILLER_37_424 ();
 sg13g2_fill_2 FILLER_37_452 ();
 sg13g2_fill_1 FILLER_37_454 ();
 sg13g2_fill_1 FILLER_37_500 ();
 sg13g2_fill_1 FILLER_37_552 ();
 sg13g2_fill_2 FILLER_37_566 ();
 sg13g2_fill_2 FILLER_37_619 ();
 sg13g2_fill_1 FILLER_37_621 ();
 sg13g2_fill_2 FILLER_37_653 ();
 sg13g2_fill_2 FILLER_37_700 ();
 sg13g2_fill_1 FILLER_37_702 ();
 sg13g2_fill_2 FILLER_37_728 ();
 sg13g2_fill_1 FILLER_37_743 ();
 sg13g2_fill_2 FILLER_37_813 ();
 sg13g2_fill_2 FILLER_37_856 ();
 sg13g2_fill_2 FILLER_37_1001 ();
 sg13g2_fill_1 FILLER_37_1003 ();
 sg13g2_fill_1 FILLER_38_8 ();
 sg13g2_fill_2 FILLER_38_18 ();
 sg13g2_fill_1 FILLER_38_20 ();
 sg13g2_fill_2 FILLER_38_57 ();
 sg13g2_fill_1 FILLER_38_59 ();
 sg13g2_fill_1 FILLER_38_78 ();
 sg13g2_fill_2 FILLER_38_97 ();
 sg13g2_fill_2 FILLER_38_107 ();
 sg13g2_fill_2 FILLER_38_116 ();
 sg13g2_fill_1 FILLER_38_118 ();
 sg13g2_fill_2 FILLER_38_146 ();
 sg13g2_fill_2 FILLER_38_185 ();
 sg13g2_fill_1 FILLER_38_187 ();
 sg13g2_fill_1 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_220 ();
 sg13g2_fill_1 FILLER_38_226 ();
 sg13g2_fill_2 FILLER_38_266 ();
 sg13g2_fill_1 FILLER_38_268 ();
 sg13g2_fill_1 FILLER_38_348 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_fill_2 FILLER_38_468 ();
 sg13g2_fill_2 FILLER_38_484 ();
 sg13g2_fill_2 FILLER_38_527 ();
 sg13g2_fill_2 FILLER_38_575 ();
 sg13g2_fill_1 FILLER_38_577 ();
 sg13g2_fill_1 FILLER_38_618 ();
 sg13g2_fill_2 FILLER_38_700 ();
 sg13g2_fill_1 FILLER_38_702 ();
 sg13g2_fill_1 FILLER_38_732 ();
 sg13g2_fill_1 FILLER_38_790 ();
 sg13g2_fill_1 FILLER_38_839 ();
 sg13g2_fill_2 FILLER_38_972 ();
 sg13g2_fill_2 FILLER_38_1001 ();
 sg13g2_fill_2 FILLER_38_1026 ();
 sg13g2_fill_1 FILLER_38_1028 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_6 ();
 sg13g2_fill_1 FILLER_39_35 ();
 sg13g2_fill_2 FILLER_39_71 ();
 sg13g2_fill_2 FILLER_39_106 ();
 sg13g2_fill_1 FILLER_39_108 ();
 sg13g2_fill_1 FILLER_39_119 ();
 sg13g2_fill_1 FILLER_39_149 ();
 sg13g2_fill_1 FILLER_39_167 ();
 sg13g2_fill_1 FILLER_39_194 ();
 sg13g2_fill_1 FILLER_39_216 ();
 sg13g2_fill_1 FILLER_39_371 ();
 sg13g2_fill_2 FILLER_39_385 ();
 sg13g2_fill_2 FILLER_39_429 ();
 sg13g2_fill_1 FILLER_39_431 ();
 sg13g2_fill_2 FILLER_39_485 ();
 sg13g2_fill_2 FILLER_39_513 ();
 sg13g2_fill_1 FILLER_39_569 ();
 sg13g2_fill_2 FILLER_39_592 ();
 sg13g2_fill_2 FILLER_39_615 ();
 sg13g2_fill_1 FILLER_39_617 ();
 sg13g2_fill_1 FILLER_39_705 ();
 sg13g2_fill_2 FILLER_39_715 ();
 sg13g2_fill_1 FILLER_39_717 ();
 sg13g2_fill_2 FILLER_39_824 ();
 sg13g2_fill_1 FILLER_39_919 ();
 sg13g2_fill_2 FILLER_39_986 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_51 ();
 sg13g2_fill_2 FILLER_40_120 ();
 sg13g2_fill_1 FILLER_40_122 ();
 sg13g2_fill_1 FILLER_40_181 ();
 sg13g2_fill_2 FILLER_40_245 ();
 sg13g2_fill_1 FILLER_40_247 ();
 sg13g2_fill_1 FILLER_40_265 ();
 sg13g2_fill_1 FILLER_40_377 ();
 sg13g2_fill_1 FILLER_40_405 ();
 sg13g2_fill_2 FILLER_40_433 ();
 sg13g2_fill_2 FILLER_40_475 ();
 sg13g2_fill_1 FILLER_40_530 ();
 sg13g2_fill_2 FILLER_40_670 ();
 sg13g2_fill_2 FILLER_40_710 ();
 sg13g2_fill_1 FILLER_40_746 ();
 sg13g2_fill_1 FILLER_40_945 ();
 sg13g2_fill_2 FILLER_40_962 ();
 sg13g2_fill_1 FILLER_40_1001 ();
 sg13g2_fill_1 FILLER_41_8 ();
 sg13g2_fill_1 FILLER_41_14 ();
 sg13g2_fill_2 FILLER_41_64 ();
 sg13g2_fill_2 FILLER_41_93 ();
 sg13g2_fill_2 FILLER_41_129 ();
 sg13g2_fill_1 FILLER_41_131 ();
 sg13g2_fill_2 FILLER_41_165 ();
 sg13g2_fill_1 FILLER_41_209 ();
 sg13g2_fill_2 FILLER_41_267 ();
 sg13g2_fill_1 FILLER_41_269 ();
 sg13g2_fill_2 FILLER_41_306 ();
 sg13g2_fill_1 FILLER_41_340 ();
 sg13g2_fill_2 FILLER_41_381 ();
 sg13g2_fill_2 FILLER_41_396 ();
 sg13g2_fill_1 FILLER_41_424 ();
 sg13g2_fill_1 FILLER_41_534 ();
 sg13g2_fill_2 FILLER_41_604 ();
 sg13g2_fill_2 FILLER_41_620 ();
 sg13g2_fill_1 FILLER_41_637 ();
 sg13g2_fill_2 FILLER_41_720 ();
 sg13g2_fill_1 FILLER_41_764 ();
 sg13g2_fill_1 FILLER_41_787 ();
 sg13g2_fill_2 FILLER_41_849 ();
 sg13g2_fill_2 FILLER_41_922 ();
 sg13g2_fill_1 FILLER_41_973 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_58 ();
 sg13g2_fill_2 FILLER_42_110 ();
 sg13g2_fill_1 FILLER_42_211 ();
 sg13g2_fill_1 FILLER_42_274 ();
 sg13g2_fill_1 FILLER_42_348 ();
 sg13g2_fill_2 FILLER_42_393 ();
 sg13g2_fill_1 FILLER_42_418 ();
 sg13g2_fill_1 FILLER_42_523 ();
 sg13g2_fill_1 FILLER_42_537 ();
 sg13g2_fill_1 FILLER_42_597 ();
 sg13g2_fill_2 FILLER_42_620 ();
 sg13g2_fill_1 FILLER_42_631 ();
 sg13g2_fill_1 FILLER_42_673 ();
 sg13g2_fill_2 FILLER_42_696 ();
 sg13g2_fill_1 FILLER_42_698 ();
 sg13g2_fill_2 FILLER_42_737 ();
 sg13g2_fill_1 FILLER_42_739 ();
 sg13g2_fill_2 FILLER_42_849 ();
 sg13g2_fill_2 FILLER_42_887 ();
 sg13g2_fill_2 FILLER_42_907 ();
 sg13g2_fill_1 FILLER_42_963 ();
 sg13g2_fill_2 FILLER_42_991 ();
 sg13g2_fill_1 FILLER_42_993 ();
 sg13g2_fill_2 FILLER_42_1027 ();
 sg13g2_fill_1 FILLER_43_4 ();
 sg13g2_fill_2 FILLER_43_66 ();
 sg13g2_fill_1 FILLER_43_68 ();
 sg13g2_fill_2 FILLER_43_99 ();
 sg13g2_fill_1 FILLER_43_101 ();
 sg13g2_fill_2 FILLER_43_107 ();
 sg13g2_fill_1 FILLER_43_109 ();
 sg13g2_fill_1 FILLER_43_120 ();
 sg13g2_fill_1 FILLER_43_134 ();
 sg13g2_fill_1 FILLER_43_140 ();
 sg13g2_fill_2 FILLER_43_155 ();
 sg13g2_fill_1 FILLER_43_157 ();
 sg13g2_fill_2 FILLER_43_172 ();
 sg13g2_fill_1 FILLER_43_183 ();
 sg13g2_fill_2 FILLER_43_232 ();
 sg13g2_fill_2 FILLER_43_275 ();
 sg13g2_fill_1 FILLER_43_277 ();
 sg13g2_fill_1 FILLER_43_342 ();
 sg13g2_fill_1 FILLER_43_359 ();
 sg13g2_fill_1 FILLER_43_393 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_fill_2 FILLER_43_446 ();
 sg13g2_fill_1 FILLER_43_507 ();
 sg13g2_fill_2 FILLER_43_529 ();
 sg13g2_fill_2 FILLER_43_559 ();
 sg13g2_fill_2 FILLER_43_588 ();
 sg13g2_fill_1 FILLER_43_590 ();
 sg13g2_fill_1 FILLER_43_610 ();
 sg13g2_fill_2 FILLER_43_634 ();
 sg13g2_fill_1 FILLER_43_659 ();
 sg13g2_fill_1 FILLER_43_721 ();
 sg13g2_fill_2 FILLER_43_740 ();
 sg13g2_fill_1 FILLER_43_816 ();
 sg13g2_fill_2 FILLER_43_884 ();
 sg13g2_fill_1 FILLER_43_886 ();
 sg13g2_fill_1 FILLER_43_946 ();
 sg13g2_fill_1 FILLER_43_1001 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_114 ();
 sg13g2_fill_1 FILLER_44_116 ();
 sg13g2_fill_2 FILLER_44_135 ();
 sg13g2_fill_2 FILLER_44_174 ();
 sg13g2_fill_1 FILLER_44_266 ();
 sg13g2_fill_1 FILLER_44_299 ();
 sg13g2_fill_1 FILLER_44_346 ();
 sg13g2_fill_1 FILLER_44_372 ();
 sg13g2_fill_2 FILLER_44_419 ();
 sg13g2_fill_2 FILLER_44_453 ();
 sg13g2_fill_1 FILLER_44_455 ();
 sg13g2_fill_2 FILLER_44_461 ();
 sg13g2_fill_1 FILLER_44_463 ();
 sg13g2_fill_1 FILLER_44_508 ();
 sg13g2_fill_2 FILLER_44_529 ();
 sg13g2_fill_2 FILLER_44_536 ();
 sg13g2_fill_1 FILLER_44_538 ();
 sg13g2_fill_2 FILLER_44_549 ();
 sg13g2_fill_1 FILLER_44_611 ();
 sg13g2_fill_1 FILLER_44_661 ();
 sg13g2_fill_2 FILLER_44_677 ();
 sg13g2_fill_2 FILLER_44_702 ();
 sg13g2_fill_1 FILLER_44_704 ();
 sg13g2_fill_1 FILLER_44_714 ();
 sg13g2_fill_2 FILLER_44_723 ();
 sg13g2_fill_1 FILLER_44_757 ();
 sg13g2_fill_1 FILLER_44_790 ();
 sg13g2_fill_2 FILLER_44_935 ();
 sg13g2_fill_2 FILLER_44_947 ();
 sg13g2_fill_2 FILLER_44_990 ();
 sg13g2_fill_1 FILLER_44_998 ();
 sg13g2_fill_2 FILLER_44_1026 ();
 sg13g2_fill_1 FILLER_44_1028 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_34 ();
 sg13g2_fill_2 FILLER_45_49 ();
 sg13g2_fill_2 FILLER_45_92 ();
 sg13g2_fill_2 FILLER_45_103 ();
 sg13g2_fill_2 FILLER_45_182 ();
 sg13g2_fill_1 FILLER_45_184 ();
 sg13g2_fill_1 FILLER_45_220 ();
 sg13g2_fill_2 FILLER_45_248 ();
 sg13g2_fill_1 FILLER_45_250 ();
 sg13g2_fill_2 FILLER_45_433 ();
 sg13g2_fill_2 FILLER_45_500 ();
 sg13g2_fill_1 FILLER_45_525 ();
 sg13g2_fill_1 FILLER_45_578 ();
 sg13g2_fill_1 FILLER_45_662 ();
 sg13g2_fill_1 FILLER_45_681 ();
 sg13g2_fill_2 FILLER_45_764 ();
 sg13g2_fill_2 FILLER_45_779 ();
 sg13g2_fill_1 FILLER_45_781 ();
 sg13g2_fill_2 FILLER_45_799 ();
 sg13g2_fill_1 FILLER_45_801 ();
 sg13g2_fill_1 FILLER_45_824 ();
 sg13g2_fill_1 FILLER_45_877 ();
 sg13g2_fill_2 FILLER_45_938 ();
 sg13g2_fill_1 FILLER_45_999 ();
 sg13g2_fill_2 FILLER_45_1023 ();
 sg13g2_fill_2 FILLER_46_8 ();
 sg13g2_fill_1 FILLER_46_10 ();
 sg13g2_fill_2 FILLER_46_23 ();
 sg13g2_fill_1 FILLER_46_52 ();
 sg13g2_fill_2 FILLER_46_134 ();
 sg13g2_fill_1 FILLER_46_163 ();
 sg13g2_fill_2 FILLER_46_199 ();
 sg13g2_fill_1 FILLER_46_248 ();
 sg13g2_fill_1 FILLER_46_276 ();
 sg13g2_fill_2 FILLER_46_309 ();
 sg13g2_fill_1 FILLER_46_348 ();
 sg13g2_fill_1 FILLER_46_380 ();
 sg13g2_fill_1 FILLER_46_399 ();
 sg13g2_fill_1 FILLER_46_486 ();
 sg13g2_fill_1 FILLER_46_496 ();
 sg13g2_fill_1 FILLER_46_502 ();
 sg13g2_fill_1 FILLER_46_529 ();
 sg13g2_fill_1 FILLER_46_534 ();
 sg13g2_fill_1 FILLER_46_591 ();
 sg13g2_fill_2 FILLER_46_722 ();
 sg13g2_fill_2 FILLER_46_760 ();
 sg13g2_fill_2 FILLER_46_780 ();
 sg13g2_fill_2 FILLER_46_810 ();
 sg13g2_fill_1 FILLER_46_812 ();
 sg13g2_fill_2 FILLER_46_855 ();
 sg13g2_fill_2 FILLER_46_925 ();
 sg13g2_fill_1 FILLER_46_971 ();
 sg13g2_fill_1 FILLER_46_984 ();
 sg13g2_fill_2 FILLER_46_1026 ();
 sg13g2_fill_1 FILLER_46_1028 ();
 sg13g2_decap_8 FILLER_47_8 ();
 sg13g2_decap_4 FILLER_47_15 ();
 sg13g2_fill_1 FILLER_47_19 ();
 sg13g2_decap_8 FILLER_47_23 ();
 sg13g2_fill_1 FILLER_47_30 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_fill_2 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_54 ();
 sg13g2_decap_8 FILLER_47_61 ();
 sg13g2_decap_8 FILLER_47_68 ();
 sg13g2_decap_4 FILLER_47_75 ();
 sg13g2_fill_2 FILLER_47_83 ();
 sg13g2_fill_1 FILLER_47_85 ();
 sg13g2_fill_2 FILLER_47_100 ();
 sg13g2_fill_1 FILLER_47_102 ();
 sg13g2_fill_1 FILLER_47_112 ();
 sg13g2_fill_2 FILLER_47_176 ();
 sg13g2_fill_2 FILLER_47_209 ();
 sg13g2_fill_2 FILLER_47_284 ();
 sg13g2_fill_1 FILLER_47_403 ();
 sg13g2_fill_2 FILLER_47_537 ();
 sg13g2_fill_2 FILLER_47_562 ();
 sg13g2_fill_1 FILLER_47_564 ();
 sg13g2_fill_1 FILLER_47_570 ();
 sg13g2_fill_2 FILLER_47_597 ();
 sg13g2_fill_1 FILLER_47_599 ();
 sg13g2_fill_2 FILLER_47_669 ();
 sg13g2_fill_1 FILLER_47_681 ();
 sg13g2_fill_1 FILLER_47_760 ();
 sg13g2_fill_1 FILLER_47_780 ();
 sg13g2_fill_1 FILLER_47_795 ();
 sg13g2_fill_1 FILLER_47_850 ();
 sg13g2_fill_1 FILLER_47_878 ();
 sg13g2_decap_8 FILLER_47_1020 ();
 sg13g2_fill_2 FILLER_47_1027 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_4 FILLER_48_77 ();
 sg13g2_fill_2 FILLER_48_81 ();
 sg13g2_decap_4 FILLER_48_87 ();
 sg13g2_fill_1 FILLER_48_91 ();
 sg13g2_fill_2 FILLER_48_121 ();
 sg13g2_fill_1 FILLER_48_123 ();
 sg13g2_fill_2 FILLER_48_182 ();
 sg13g2_fill_1 FILLER_48_292 ();
 sg13g2_fill_2 FILLER_48_320 ();
 sg13g2_fill_1 FILLER_48_351 ();
 sg13g2_fill_1 FILLER_48_367 ();
 sg13g2_fill_1 FILLER_48_394 ();
 sg13g2_fill_1 FILLER_48_422 ();
 sg13g2_fill_1 FILLER_48_451 ();
 sg13g2_fill_1 FILLER_48_484 ();
 sg13g2_fill_1 FILLER_48_519 ();
 sg13g2_fill_2 FILLER_48_537 ();
 sg13g2_fill_2 FILLER_48_573 ();
 sg13g2_fill_1 FILLER_48_647 ();
 sg13g2_fill_1 FILLER_48_661 ();
 sg13g2_fill_2 FILLER_48_667 ();
 sg13g2_fill_1 FILLER_48_669 ();
 sg13g2_fill_2 FILLER_48_697 ();
 sg13g2_fill_1 FILLER_48_699 ();
 sg13g2_fill_1 FILLER_48_728 ();
 sg13g2_fill_2 FILLER_48_738 ();
 sg13g2_fill_1 FILLER_48_740 ();
 sg13g2_fill_2 FILLER_48_768 ();
 sg13g2_fill_1 FILLER_48_770 ();
 sg13g2_fill_2 FILLER_48_934 ();
 sg13g2_decap_8 FILLER_48_1007 ();
 sg13g2_decap_8 FILLER_48_1014 ();
 sg13g2_decap_8 FILLER_48_1021 ();
 sg13g2_fill_1 FILLER_48_1028 ();
 sg13g2_decap_8 FILLER_49_5 ();
 sg13g2_decap_8 FILLER_49_12 ();
 sg13g2_decap_8 FILLER_49_19 ();
 sg13g2_decap_8 FILLER_49_26 ();
 sg13g2_decap_8 FILLER_49_33 ();
 sg13g2_decap_8 FILLER_49_40 ();
 sg13g2_decap_8 FILLER_49_47 ();
 sg13g2_decap_8 FILLER_49_54 ();
 sg13g2_decap_8 FILLER_49_61 ();
 sg13g2_decap_8 FILLER_49_68 ();
 sg13g2_decap_8 FILLER_49_75 ();
 sg13g2_decap_8 FILLER_49_82 ();
 sg13g2_decap_8 FILLER_49_89 ();
 sg13g2_fill_2 FILLER_49_96 ();
 sg13g2_fill_1 FILLER_49_98 ();
 sg13g2_fill_2 FILLER_49_369 ();
 sg13g2_fill_2 FILLER_49_397 ();
 sg13g2_fill_2 FILLER_49_421 ();
 sg13g2_fill_1 FILLER_49_423 ();
 sg13g2_fill_2 FILLER_49_464 ();
 sg13g2_fill_1 FILLER_49_466 ();
 sg13g2_fill_1 FILLER_49_500 ();
 sg13g2_fill_2 FILLER_49_555 ();
 sg13g2_fill_2 FILLER_49_620 ();
 sg13g2_fill_1 FILLER_49_622 ();
 sg13g2_fill_2 FILLER_49_660 ();
 sg13g2_fill_2 FILLER_49_672 ();
 sg13g2_fill_1 FILLER_49_674 ();
 sg13g2_fill_2 FILLER_49_680 ();
 sg13g2_fill_2 FILLER_49_707 ();
 sg13g2_fill_1 FILLER_49_709 ();
 sg13g2_fill_2 FILLER_49_750 ();
 sg13g2_fill_1 FILLER_49_752 ();
 sg13g2_fill_1 FILLER_49_894 ();
 sg13g2_fill_1 FILLER_49_924 ();
 sg13g2_fill_2 FILLER_49_943 ();
 sg13g2_decap_8 FILLER_49_1000 ();
 sg13g2_decap_8 FILLER_49_1007 ();
 sg13g2_decap_8 FILLER_49_1014 ();
 sg13g2_decap_8 FILLER_49_1021 ();
 sg13g2_fill_1 FILLER_49_1028 ();
 assign uio_oe[0] = net24;
 assign uio_oe[1] = net25;
 assign uio_oe[2] = net26;
 assign uio_oe[3] = net27;
 assign uio_oe[4] = net28;
 assign uio_oe[5] = net29;
 assign uio_oe[6] = net30;
 assign uio_oe[7] = net757;
 assign uio_out[0] = net31;
 assign uio_out[1] = net32;
 assign uio_out[2] = net33;
 assign uio_out[3] = net34;
 assign uio_out[4] = net35;
 assign uio_out[5] = net36;
 assign uio_out[6] = net37;
 assign uo_out[2] = net38;
 assign uo_out[6] = net39;
endmodule
